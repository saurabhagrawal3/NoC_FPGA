//---------------------------------------------------------------------------------------
// uart transmit module  
//
//---------------------------------------------------------------------------------------

module uart_tx  
(
	clock, reset,
	ce_32, tx_data, new_tx_data, 
	ser_out, tx_busy
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
input			ce_32;			// baud rate multiplyed by 16 - generated by baud module 
input	[15:0]	tx_data;		// data byte to transmit 
input			new_tx_data;	// asserted to indicate that there is a new data byte for transmission 
output			ser_out;		// serial data output 
output 			tx_busy;		// signs that transmitter is busy 

// internal wires 
wire ce_1;		// clock enable at bit rate 

// internal registers 
reg ser_out;
reg tx_busy;
reg [4:0]	count32;
reg [4:0]	bit_count;
reg [16:0]	data_buf;
reg reg_new_tx_data;
//---------------------------------------------------------------------------------------
// module implementation 
// a counter to count 16 pulses of ce_32 to generate the ce_1 pulse 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		count32 <= 5'b0;
	else if (tx_busy & ce_32)
		count32 <= count32 + 5'b1;
	else if (~tx_busy)
		count32 <= 5'b0;
end 

// ce_1 pulse indicating output data bit should be updated 
assign ce_1 = (count32 == 5'b11111) & ce_32;

// tx_busy flag 
always @ (posedge clock)
begin
	reg_new_tx_data <= new_tx_data;
	if (reset) 
		tx_busy <= 1'b0;
	else if (~tx_busy & new_tx_data)
		tx_busy <= 1'b1;
	else if (tx_busy & (bit_count == 17) & ce_1)
		tx_busy <= 1'b0;
end 

// output bit counter 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		bit_count <= 5'h0;
	else if (tx_busy & ce_1)
		bit_count <= bit_count + 5'h1;
	else if (~tx_busy) 
		bit_count <= 5'h0;
end 

// data shift register 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		data_buf <= 17'b0;
	else if (~tx_busy & new_tx_data)//(~(tx_busy | new_tx_data))
		data_buf <= {tx_data, 1'b0};
	else if (tx_busy & ce_1)
		data_buf <= {1'b1, data_buf[16:1]};
end 

// output data bit 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		ser_out <= 1'b1;
	else if (tx_busy)
		ser_out <= data_buf[0];
	else 
		ser_out <= 1'b1;
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------
