`timescale 1ns / 1ps


`include "connect_parameters.v"
`include "matrix_vector_mult_parameters.v"


module mult_top_64(
   reset,
   clk,
   max_iteration,
   data_in,
   data_o,
   done
  );
  
  
  localparam RAM_ADDR_BITS= `RAM_ADDR_BITS; 
  localparam RAM_WIDTH = `RAM_WIDTH; 
  localparam VECTOR_SIZE = `VECTOR_SIZE;
  localparam folding_factor = `FOLDING_FACTOR;
  localparam vertex_width = `VERTEX_WIDTH;
  localparam vc_bits = 1;//(`NUM_VCS > 1) ? $clog2(`NUM_VCS) : 1;
  localparam dest_bits = `ADDR_WIDTH;//$clog2(`NUM_USER_RECV_PORTS);
  localparam flit_port_width = 2 /*valid and tail bits*/+ `FLIT_DATA_WIDTH + dest_bits + vc_bits;
   
  input clk, reset;
  input [VECTOR_SIZE-1:0] data_in;
  input [15:0] max_iteration;
  output [VECTOR_SIZE-1:0] data_o;
  output done;
  
  wire rst_n;
  
  assign rst_n = !reset;
  
  
 wire [flit_port_width-1:0]  send_ports_0_putFlit_flit_in,  send_ports_1_putFlit_flit_in,  send_ports_2_putFlit_flit_in,  send_ports_3_putFlit_flit_in,  send_ports_4_putFlit_flit_in,  send_ports_5_putFlit_flit_in,  send_ports_6_putFlit_flit_in,  send_ports_7_putFlit_flit_in,  send_ports_8_putFlit_flit_in,  send_ports_9_putFlit_flit_in,  send_ports_10_putFlit_flit_in,  send_ports_11_putFlit_flit_in,  send_ports_12_putFlit_flit_in,  send_ports_13_putFlit_flit_in,  send_ports_14_putFlit_flit_in,  send_ports_15_putFlit_flit_in,  send_ports_16_putFlit_flit_in,  send_ports_17_putFlit_flit_in,  send_ports_18_putFlit_flit_in,  send_ports_19_putFlit_flit_in,  send_ports_20_putFlit_flit_in,  send_ports_21_putFlit_flit_in,  send_ports_22_putFlit_flit_in,  send_ports_23_putFlit_flit_in,  send_ports_24_putFlit_flit_in,  send_ports_25_putFlit_flit_in,  send_ports_26_putFlit_flit_in,  send_ports_27_putFlit_flit_in,  send_ports_28_putFlit_flit_in,  send_ports_29_putFlit_flit_in,  send_ports_30_putFlit_flit_in,  send_ports_31_putFlit_flit_in,  send_ports_32_putFlit_flit_in,  send_ports_33_putFlit_flit_in,  send_ports_34_putFlit_flit_in,  send_ports_35_putFlit_flit_in,  send_ports_36_putFlit_flit_in,  send_ports_37_putFlit_flit_in,  send_ports_38_putFlit_flit_in,  send_ports_39_putFlit_flit_in,  send_ports_40_putFlit_flit_in,  send_ports_41_putFlit_flit_in,  send_ports_42_putFlit_flit_in,  send_ports_43_putFlit_flit_in,  send_ports_44_putFlit_flit_in,  send_ports_45_putFlit_flit_in,  send_ports_46_putFlit_flit_in,  send_ports_47_putFlit_flit_in,  send_ports_48_putFlit_flit_in,  send_ports_49_putFlit_flit_in,  send_ports_50_putFlit_flit_in,  send_ports_51_putFlit_flit_in,  send_ports_52_putFlit_flit_in,  send_ports_53_putFlit_flit_in,  send_ports_54_putFlit_flit_in,  send_ports_55_putFlit_flit_in,  send_ports_56_putFlit_flit_in,  send_ports_57_putFlit_flit_in,  send_ports_58_putFlit_flit_in,  send_ports_59_putFlit_flit_in,  send_ports_60_putFlit_flit_in,  send_ports_61_putFlit_flit_in,  send_ports_62_putFlit_flit_in,  send_ports_63_putFlit_flit_in;
  
  
wire  EN_send_ports_0_putFlit,  EN_send_ports_1_putFlit,  EN_send_ports_2_putFlit,  EN_send_ports_3_putFlit,  EN_send_ports_4_putFlit,  EN_send_ports_5_putFlit,  EN_send_ports_6_putFlit,  EN_send_ports_7_putFlit,  EN_send_ports_8_putFlit,  EN_send_ports_9_putFlit,  EN_send_ports_10_putFlit,  EN_send_ports_11_putFlit,  EN_send_ports_12_putFlit,  EN_send_ports_13_putFlit,  EN_send_ports_14_putFlit,  EN_send_ports_15_putFlit,  EN_send_ports_16_putFlit,  EN_send_ports_17_putFlit,  EN_send_ports_18_putFlit,  EN_send_ports_19_putFlit,  EN_send_ports_20_putFlit,  EN_send_ports_21_putFlit,  EN_send_ports_22_putFlit,  EN_send_ports_23_putFlit,  EN_send_ports_24_putFlit,  EN_send_ports_25_putFlit,  EN_send_ports_26_putFlit,  EN_send_ports_27_putFlit,  EN_send_ports_28_putFlit,  EN_send_ports_29_putFlit,  EN_send_ports_30_putFlit,  EN_send_ports_31_putFlit,  EN_send_ports_32_putFlit,  EN_send_ports_33_putFlit,  EN_send_ports_34_putFlit,  EN_send_ports_35_putFlit,  EN_send_ports_36_putFlit,  EN_send_ports_37_putFlit,  EN_send_ports_38_putFlit,  EN_send_ports_39_putFlit,  EN_send_ports_40_putFlit,  EN_send_ports_41_putFlit,  EN_send_ports_42_putFlit,  EN_send_ports_43_putFlit,  EN_send_ports_44_putFlit,  EN_send_ports_45_putFlit,  EN_send_ports_46_putFlit,  EN_send_ports_47_putFlit,  EN_send_ports_48_putFlit,  EN_send_ports_49_putFlit,  EN_send_ports_50_putFlit,  EN_send_ports_51_putFlit,  EN_send_ports_52_putFlit,  EN_send_ports_53_putFlit,  EN_send_ports_54_putFlit,  EN_send_ports_55_putFlit,  EN_send_ports_56_putFlit,  EN_send_ports_57_putFlit,  EN_send_ports_58_putFlit,  EN_send_ports_59_putFlit,  EN_send_ports_60_putFlit,  EN_send_ports_61_putFlit,  EN_send_ports_62_putFlit,  EN_send_ports_63_putFlit; 


wire [1:0]  send_ports_0_getNonFullVCs,  send_ports_1_getNonFullVCs,  send_ports_2_getNonFullVCs,  send_ports_3_getNonFullVCs,  send_ports_4_getNonFullVCs,  send_ports_5_getNonFullVCs,  send_ports_6_getNonFullVCs,  send_ports_7_getNonFullVCs,  send_ports_8_getNonFullVCs,  send_ports_9_getNonFullVCs,  send_ports_10_getNonFullVCs,  send_ports_11_getNonFullVCs,  send_ports_12_getNonFullVCs,  send_ports_13_getNonFullVCs,  send_ports_14_getNonFullVCs,  send_ports_15_getNonFullVCs,  send_ports_16_getNonFullVCs,  send_ports_17_getNonFullVCs,  send_ports_18_getNonFullVCs,  send_ports_19_getNonFullVCs,  send_ports_20_getNonFullVCs,  send_ports_21_getNonFullVCs,  send_ports_22_getNonFullVCs,  send_ports_23_getNonFullVCs,  send_ports_24_getNonFullVCs,  send_ports_25_getNonFullVCs,  send_ports_26_getNonFullVCs,  send_ports_27_getNonFullVCs,  send_ports_28_getNonFullVCs,  send_ports_29_getNonFullVCs,  send_ports_30_getNonFullVCs,  send_ports_31_getNonFullVCs,  send_ports_32_getNonFullVCs,  send_ports_33_getNonFullVCs,  send_ports_34_getNonFullVCs,  send_ports_35_getNonFullVCs,  send_ports_36_getNonFullVCs,  send_ports_37_getNonFullVCs,  send_ports_38_getNonFullVCs,  send_ports_39_getNonFullVCs,  send_ports_40_getNonFullVCs,  send_ports_41_getNonFullVCs,  send_ports_42_getNonFullVCs,  send_ports_43_getNonFullVCs,  send_ports_44_getNonFullVCs,  send_ports_45_getNonFullVCs,  send_ports_46_getNonFullVCs,  send_ports_47_getNonFullVCs,  send_ports_48_getNonFullVCs,  send_ports_49_getNonFullVCs,  send_ports_50_getNonFullVCs,  send_ports_51_getNonFullVCs,  send_ports_52_getNonFullVCs,  send_ports_53_getNonFullVCs,  send_ports_54_getNonFullVCs,  send_ports_55_getNonFullVCs,  send_ports_56_getNonFullVCs,  send_ports_57_getNonFullVCs,  send_ports_58_getNonFullVCs,  send_ports_59_getNonFullVCs,  send_ports_60_getNonFullVCs,  send_ports_61_getNonFullVCs,  send_ports_62_getNonFullVCs,  send_ports_63_getNonFullVCs;

wire [flit_port_width-1:0]  recv_ports_0_getFlit,  recv_ports_1_getFlit,  recv_ports_2_getFlit,  recv_ports_3_getFlit,  recv_ports_4_getFlit,  recv_ports_5_getFlit,  recv_ports_6_getFlit,  recv_ports_7_getFlit,  recv_ports_8_getFlit,  recv_ports_9_getFlit,  recv_ports_10_getFlit,  recv_ports_11_getFlit,  recv_ports_12_getFlit,  recv_ports_13_getFlit,  recv_ports_14_getFlit,  recv_ports_15_getFlit,  recv_ports_16_getFlit,  recv_ports_17_getFlit,  recv_ports_18_getFlit,  recv_ports_19_getFlit,  recv_ports_20_getFlit,  recv_ports_21_getFlit,  recv_ports_22_getFlit,  recv_ports_23_getFlit,  recv_ports_24_getFlit,  recv_ports_25_getFlit,  recv_ports_26_getFlit,  recv_ports_27_getFlit,  recv_ports_28_getFlit,  recv_ports_29_getFlit,  recv_ports_30_getFlit,  recv_ports_31_getFlit,  recv_ports_32_getFlit,  recv_ports_33_getFlit,  recv_ports_34_getFlit,  recv_ports_35_getFlit,  recv_ports_36_getFlit,  recv_ports_37_getFlit,  recv_ports_38_getFlit,  recv_ports_39_getFlit,  recv_ports_40_getFlit,  recv_ports_41_getFlit,  recv_ports_42_getFlit,  recv_ports_43_getFlit,  recv_ports_44_getFlit,  recv_ports_45_getFlit,  recv_ports_46_getFlit,  recv_ports_47_getFlit,  recv_ports_48_getFlit,  recv_ports_49_getFlit,  recv_ports_50_getFlit,  recv_ports_51_getFlit,  recv_ports_52_getFlit,  recv_ports_53_getFlit,  recv_ports_54_getFlit,  recv_ports_55_getFlit,  recv_ports_56_getFlit,  recv_ports_57_getFlit,  recv_ports_58_getFlit,  recv_ports_59_getFlit,  recv_ports_60_getFlit,  recv_ports_61_getFlit,  recv_ports_62_getFlit,  recv_ports_63_getFlit;

wire [dest_bits-1:0] recv_ports_info_0_getRecvPortID, recv_ports_info_1_getRecvPortID, recv_ports_info_2_getRecvPortID, recv_ports_info_3_getRecvPortID, recv_ports_info_4_getRecvPortID, recv_ports_info_5_getRecvPortID, recv_ports_info_6_getRecvPortID, recv_ports_info_7_getRecvPortID, recv_ports_info_8_getRecvPortID, recv_ports_info_9_getRecvPortID, recv_ports_info_10_getRecvPortID, recv_ports_info_11_getRecvPortID, recv_ports_info_12_getRecvPortID, recv_ports_info_13_getRecvPortID, recv_ports_info_14_getRecvPortID, recv_ports_info_15_getRecvPortID, recv_ports_info_16_getRecvPortID, recv_ports_info_17_getRecvPortID, recv_ports_info_18_getRecvPortID, recv_ports_info_19_getRecvPortID, recv_ports_info_20_getRecvPortID, recv_ports_info_21_getRecvPortID, recv_ports_info_22_getRecvPortID, recv_ports_info_23_getRecvPortID, recv_ports_info_24_getRecvPortID, recv_ports_info_25_getRecvPortID, recv_ports_info_26_getRecvPortID, recv_ports_info_27_getRecvPortID, recv_ports_info_28_getRecvPortID, recv_ports_info_29_getRecvPortID, recv_ports_info_30_getRecvPortID, recv_ports_info_31_getRecvPortID, recv_ports_info_32_getRecvPortID, recv_ports_info_33_getRecvPortID, recv_ports_info_34_getRecvPortID, recv_ports_info_35_getRecvPortID, recv_ports_info_36_getRecvPortID, recv_ports_info_37_getRecvPortID, recv_ports_info_38_getRecvPortID, recv_ports_info_39_getRecvPortID, recv_ports_info_40_getRecvPortID, recv_ports_info_41_getRecvPortID, recv_ports_info_42_getRecvPortID, recv_ports_info_43_getRecvPortID, recv_ports_info_44_getRecvPortID, recv_ports_info_45_getRecvPortID, recv_ports_info_46_getRecvPortID, recv_ports_info_47_getRecvPortID, recv_ports_info_48_getRecvPortID, recv_ports_info_49_getRecvPortID, recv_ports_info_50_getRecvPortID, recv_ports_info_51_getRecvPortID, recv_ports_info_52_getRecvPortID, recv_ports_info_53_getRecvPortID, recv_ports_info_54_getRecvPortID, recv_ports_info_55_getRecvPortID, recv_ports_info_56_getRecvPortID, recv_ports_info_57_getRecvPortID, recv_ports_info_58_getRecvPortID, recv_ports_info_59_getRecvPortID, recv_ports_info_60_getRecvPortID, recv_ports_info_61_getRecvPortID, recv_ports_info_62_getRecvPortID, recv_ports_info_63_getRecvPortID;


wire  EN_recv_ports_0_getFlit,  EN_recv_ports_1_getFlit,  EN_recv_ports_2_getFlit,  EN_recv_ports_3_getFlit,  EN_recv_ports_4_getFlit,  EN_recv_ports_5_getFlit,  EN_recv_ports_6_getFlit,  EN_recv_ports_7_getFlit,  EN_recv_ports_8_getFlit,  EN_recv_ports_9_getFlit,  EN_recv_ports_10_getFlit,  EN_recv_ports_11_getFlit,  EN_recv_ports_12_getFlit,  EN_recv_ports_13_getFlit,  EN_recv_ports_14_getFlit,  EN_recv_ports_15_getFlit,  EN_recv_ports_16_getFlit,  EN_recv_ports_17_getFlit,  EN_recv_ports_18_getFlit,  EN_recv_ports_19_getFlit,  EN_recv_ports_20_getFlit,  EN_recv_ports_21_getFlit,  EN_recv_ports_22_getFlit,  EN_recv_ports_23_getFlit,  EN_recv_ports_24_getFlit,  EN_recv_ports_25_getFlit,  EN_recv_ports_26_getFlit,  EN_recv_ports_27_getFlit,  EN_recv_ports_28_getFlit,  EN_recv_ports_29_getFlit,  EN_recv_ports_30_getFlit,  EN_recv_ports_31_getFlit,  EN_recv_ports_32_getFlit,  EN_recv_ports_33_getFlit,  EN_recv_ports_34_getFlit,  EN_recv_ports_35_getFlit,  EN_recv_ports_36_getFlit,  EN_recv_ports_37_getFlit,  EN_recv_ports_38_getFlit,  EN_recv_ports_39_getFlit,  EN_recv_ports_40_getFlit,  EN_recv_ports_41_getFlit,  EN_recv_ports_42_getFlit,  EN_recv_ports_43_getFlit,  EN_recv_ports_44_getFlit,  EN_recv_ports_45_getFlit,  EN_recv_ports_46_getFlit,  EN_recv_ports_47_getFlit,  EN_recv_ports_48_getFlit,  EN_recv_ports_49_getFlit,  EN_recv_ports_50_getFlit,  EN_recv_ports_51_getFlit,  EN_recv_ports_52_getFlit,  EN_recv_ports_53_getFlit,  EN_recv_ports_54_getFlit,  EN_recv_ports_55_getFlit,  EN_recv_ports_56_getFlit,  EN_recv_ports_57_getFlit,  EN_recv_ports_58_getFlit,  EN_recv_ports_59_getFlit,  EN_recv_ports_60_getFlit,  EN_recv_ports_61_getFlit,  EN_recv_ports_62_getFlit,  EN_recv_ports_63_getFlit;

wire [RAM_ADDR_BITS-1:0] LUT_address_0, LUT_address_1, LUT_address_2, LUT_address_3, LUT_address_4, LUT_address_5, LUT_address_6, LUT_address_7, LUT_address_8, LUT_address_9, LUT_address_10, LUT_address_11, LUT_address_12, LUT_address_13, LUT_address_14, LUT_address_15, LUT_address_16, LUT_address_17, LUT_address_18, LUT_address_19, LUT_address_20, LUT_address_21, LUT_address_22, LUT_address_23, LUT_address_24, LUT_address_25, LUT_address_26, LUT_address_27, LUT_address_28, LUT_address_29, LUT_address_30, LUT_address_31, LUT_address_32, LUT_address_33, LUT_address_34, LUT_address_35, LUT_address_36, LUT_address_37, LUT_address_38, LUT_address_39, LUT_address_40, LUT_address_41, LUT_address_42, LUT_address_43, LUT_address_44, LUT_address_45, LUT_address_46, LUT_address_47, LUT_address_48, LUT_address_49, LUT_address_50, LUT_address_51, LUT_address_52, LUT_address_53, LUT_address_54, LUT_address_55, LUT_address_56, LUT_address_57, LUT_address_58, LUT_address_59, LUT_address_60, LUT_address_61, LUT_address_62, LUT_address_63;

wire [RAM_WIDTH-1:0] LUT_output_data_0, LUT_output_data_1, LUT_output_data_2, LUT_output_data_3, LUT_output_data_4, LUT_output_data_5, LUT_output_data_6, LUT_output_data_7, LUT_output_data_8, LUT_output_data_9, LUT_output_data_10, LUT_output_data_11, LUT_output_data_12, LUT_output_data_13, LUT_output_data_14, LUT_output_data_15, LUT_output_data_16, LUT_output_data_17, LUT_output_data_18, LUT_output_data_19, LUT_output_data_20, LUT_output_data_21, LUT_output_data_22, LUT_output_data_23, LUT_output_data_24, LUT_output_data_25, LUT_output_data_26, LUT_output_data_27, LUT_output_data_28, LUT_output_data_29, LUT_output_data_30, LUT_output_data_31, LUT_output_data_32, LUT_output_data_33, LUT_output_data_34, LUT_output_data_35, LUT_output_data_36, LUT_output_data_37, LUT_output_data_38, LUT_output_data_39, LUT_output_data_40, LUT_output_data_41, LUT_output_data_42, LUT_output_data_43, LUT_output_data_44, LUT_output_data_45, LUT_output_data_46, LUT_output_data_47, LUT_output_data_48, LUT_output_data_49, LUT_output_data_50, LUT_output_data_51, LUT_output_data_52, LUT_output_data_53, LUT_output_data_54, LUT_output_data_55, LUT_output_data_56, LUT_output_data_57, LUT_output_data_58, LUT_output_data_59, LUT_output_data_60, LUT_output_data_61, LUT_output_data_62, LUT_output_data_63;

wire [folding_factor*vertex_width - 1:0] vertex_63, vertex_62, vertex_61, vertex_60, vertex_59, vertex_58, vertex_57, vertex_56, vertex_55, vertex_54, vertex_53, vertex_52, vertex_51, vertex_50, vertex_49, vertex_48, vertex_47, vertex_46, vertex_45, vertex_44, vertex_43, vertex_42, vertex_41, vertex_40, vertex_39, vertex_38, vertex_37, vertex_36, vertex_35, vertex_34, vertex_33, vertex_32, vertex_31, vertex_30, vertex_29, vertex_28, vertex_27, vertex_26, vertex_25, vertex_24, vertex_23, vertex_22, vertex_21, vertex_20, vertex_19, vertex_18, vertex_17, vertex_16, vertex_15, vertex_14, vertex_13, vertex_12, vertex_11, vertex_10, vertex_9, vertex_8, vertex_7, vertex_6, vertex_5, vertex_4, vertex_3, vertex_2, vertex_1, vertex_0;


wire [folding_factor*vertex_width - 1:0] getVertex_0, getVertex_1, getVertex_2, getVertex_3, getVertex_4, getVertex_5, getVertex_6, getVertex_7, getVertex_8, getVertex_9, getVertex_10, getVertex_11, getVertex_12, getVertex_13, getVertex_14, getVertex_15, getVertex_16, getVertex_17, getVertex_18, getVertex_19, getVertex_20, getVertex_21, getVertex_22, getVertex_23, getVertex_24, getVertex_25, getVertex_26, getVertex_27, getVertex_28, getVertex_29, getVertex_30, getVertex_31, getVertex_32, getVertex_33, getVertex_34, getVertex_35, getVertex_36, getVertex_37, getVertex_38, getVertex_39, getVertex_40, getVertex_41, getVertex_42, getVertex_43, getVertex_44, getVertex_45, getVertex_46, getVertex_47, getVertex_48, getVertex_49, getVertex_50, getVertex_51, getVertex_52, getVertex_53, getVertex_54, getVertex_55, getVertex_56, getVertex_57, getVertex_58, getVertex_59, getVertex_60, getVertex_61, getVertex_62, getVertex_63;


genvar i;
generate
for (i=0; i<folding_factor; i=i+1) 
  begin:m
	assign data_o[(folding_factor-i)*vertex_width*64-1:(folding_factor-i-1)*vertex_width*64] = {vertex_0[(i+1)*vertex_width-1:i*vertex_width], vertex_1[(i+1)*vertex_width-1:i*vertex_width], vertex_2[(i+1)*vertex_width-1:i*vertex_width], vertex_3[(i+1)*vertex_width-1:i*vertex_width], vertex_4[(i+1)*vertex_width-1:i*vertex_width], vertex_5[(i+1)*vertex_width-1:i*vertex_width], vertex_6[(i+1)*vertex_width-1:i*vertex_width], vertex_7[(i+1)*vertex_width-1:i*vertex_width], vertex_8[(i+1)*vertex_width-1:i*vertex_width], vertex_9[(i+1)*vertex_width-1:i*vertex_width], vertex_10[(i+1)*vertex_width-1:i*vertex_width], vertex_11[(i+1)*vertex_width-1:i*vertex_width], vertex_12[(i+1)*vertex_width-1:i*vertex_width], vertex_13[(i+1)*vertex_width-1:i*vertex_width], vertex_14[(i+1)*vertex_width-1:i*vertex_width], vertex_15[(i+1)*vertex_width-1:i*vertex_width], vertex_16[(i+1)*vertex_width-1:i*vertex_width], vertex_17[(i+1)*vertex_width-1:i*vertex_width], vertex_18[(i+1)*vertex_width-1:i*vertex_width], vertex_19[(i+1)*vertex_width-1:i*vertex_width], vertex_20[(i+1)*vertex_width-1:i*vertex_width], vertex_21[(i+1)*vertex_width-1:i*vertex_width], vertex_22[(i+1)*vertex_width-1:i*vertex_width], vertex_23[(i+1)*vertex_width-1:i*vertex_width], vertex_24[(i+1)*vertex_width-1:i*vertex_width], vertex_25[(i+1)*vertex_width-1:i*vertex_width], vertex_26[(i+1)*vertex_width-1:i*vertex_width], vertex_27[(i+1)*vertex_width-1:i*vertex_width], vertex_28[(i+1)*vertex_width-1:i*vertex_width], vertex_29[(i+1)*vertex_width-1:i*vertex_width], vertex_30[(i+1)*vertex_width-1:i*vertex_width], vertex_31[(i+1)*vertex_width-1:i*vertex_width], vertex_32[(i+1)*vertex_width-1:i*vertex_width], vertex_33[(i+1)*vertex_width-1:i*vertex_width], vertex_34[(i+1)*vertex_width-1:i*vertex_width], vertex_35[(i+1)*vertex_width-1:i*vertex_width], vertex_36[(i+1)*vertex_width-1:i*vertex_width], vertex_37[(i+1)*vertex_width-1:i*vertex_width], vertex_38[(i+1)*vertex_width-1:i*vertex_width], vertex_39[(i+1)*vertex_width-1:i*vertex_width], vertex_40[(i+1)*vertex_width-1:i*vertex_width], vertex_41[(i+1)*vertex_width-1:i*vertex_width], vertex_42[(i+1)*vertex_width-1:i*vertex_width], vertex_43[(i+1)*vertex_width-1:i*vertex_width], vertex_44[(i+1)*vertex_width-1:i*vertex_width], vertex_45[(i+1)*vertex_width-1:i*vertex_width], vertex_46[(i+1)*vertex_width-1:i*vertex_width], vertex_47[(i+1)*vertex_width-1:i*vertex_width], vertex_48[(i+1)*vertex_width-1:i*vertex_width], vertex_49[(i+1)*vertex_width-1:i*vertex_width], vertex_50[(i+1)*vertex_width-1:i*vertex_width], vertex_51[(i+1)*vertex_width-1:i*vertex_width], vertex_52[(i+1)*vertex_width-1:i*vertex_width], vertex_53[(i+1)*vertex_width-1:i*vertex_width], vertex_54[(i+1)*vertex_width-1:i*vertex_width], vertex_55[(i+1)*vertex_width-1:i*vertex_width], vertex_56[(i+1)*vertex_width-1:i*vertex_width], vertex_57[(i+1)*vertex_width-1:i*vertex_width], vertex_58[(i+1)*vertex_width-1:i*vertex_width], vertex_59[(i+1)*vertex_width-1:i*vertex_width], vertex_60[(i+1)*vertex_width-1:i*vertex_width], vertex_61[(i+1)*vertex_width-1:i*vertex_width], vertex_62[(i+1)*vertex_width-1:i*vertex_width], vertex_63[(i+1)*vertex_width-1:i*vertex_width]};

	assign {getVertex_0[(i+1)*vertex_width-1:i*vertex_width], getVertex_1[(i+1)*vertex_width-1:i*vertex_width], getVertex_2[(i+1)*vertex_width-1:i*vertex_width], getVertex_3[(i+1)*vertex_width-1:i*vertex_width], getVertex_4[(i+1)*vertex_width-1:i*vertex_width], getVertex_5[(i+1)*vertex_width-1:i*vertex_width], getVertex_6[(i+1)*vertex_width-1:i*vertex_width], getVertex_7[(i+1)*vertex_width-1:i*vertex_width], getVertex_8[(i+1)*vertex_width-1:i*vertex_width], getVertex_9[(i+1)*vertex_width-1:i*vertex_width], getVertex_10[(i+1)*vertex_width-1:i*vertex_width], getVertex_11[(i+1)*vertex_width-1:i*vertex_width], getVertex_12[(i+1)*vertex_width-1:i*vertex_width], getVertex_13[(i+1)*vertex_width-1:i*vertex_width], getVertex_14[(i+1)*vertex_width-1:i*vertex_width], getVertex_15[(i+1)*vertex_width-1:i*vertex_width], getVertex_16[(i+1)*vertex_width-1:i*vertex_width], getVertex_17[(i+1)*vertex_width-1:i*vertex_width], getVertex_18[(i+1)*vertex_width-1:i*vertex_width], getVertex_19[(i+1)*vertex_width-1:i*vertex_width], getVertex_20[(i+1)*vertex_width-1:i*vertex_width], getVertex_21[(i+1)*vertex_width-1:i*vertex_width], getVertex_22[(i+1)*vertex_width-1:i*vertex_width], getVertex_23[(i+1)*vertex_width-1:i*vertex_width], getVertex_24[(i+1)*vertex_width-1:i*vertex_width], getVertex_25[(i+1)*vertex_width-1:i*vertex_width], getVertex_26[(i+1)*vertex_width-1:i*vertex_width], getVertex_27[(i+1)*vertex_width-1:i*vertex_width], getVertex_28[(i+1)*vertex_width-1:i*vertex_width], getVertex_29[(i+1)*vertex_width-1:i*vertex_width], getVertex_30[(i+1)*vertex_width-1:i*vertex_width], getVertex_31[(i+1)*vertex_width-1:i*vertex_width], getVertex_32[(i+1)*vertex_width-1:i*vertex_width], getVertex_33[(i+1)*vertex_width-1:i*vertex_width], getVertex_34[(i+1)*vertex_width-1:i*vertex_width], getVertex_35[(i+1)*vertex_width-1:i*vertex_width], getVertex_36[(i+1)*vertex_width-1:i*vertex_width], getVertex_37[(i+1)*vertex_width-1:i*vertex_width], getVertex_38[(i+1)*vertex_width-1:i*vertex_width], getVertex_39[(i+1)*vertex_width-1:i*vertex_width], getVertex_40[(i+1)*vertex_width-1:i*vertex_width], getVertex_41[(i+1)*vertex_width-1:i*vertex_width], getVertex_42[(i+1)*vertex_width-1:i*vertex_width], getVertex_43[(i+1)*vertex_width-1:i*vertex_width], getVertex_44[(i+1)*vertex_width-1:i*vertex_width], getVertex_45[(i+1)*vertex_width-1:i*vertex_width], getVertex_46[(i+1)*vertex_width-1:i*vertex_width], getVertex_47[(i+1)*vertex_width-1:i*vertex_width], getVertex_48[(i+1)*vertex_width-1:i*vertex_width], getVertex_49[(i+1)*vertex_width-1:i*vertex_width], getVertex_50[(i+1)*vertex_width-1:i*vertex_width], getVertex_51[(i+1)*vertex_width-1:i*vertex_width], getVertex_52[(i+1)*vertex_width-1:i*vertex_width], getVertex_53[(i+1)*vertex_width-1:i*vertex_width], getVertex_54[(i+1)*vertex_width-1:i*vertex_width], getVertex_55[(i+1)*vertex_width-1:i*vertex_width], getVertex_56[(i+1)*vertex_width-1:i*vertex_width], getVertex_57[(i+1)*vertex_width-1:i*vertex_width], getVertex_58[(i+1)*vertex_width-1:i*vertex_width], getVertex_59[(i+1)*vertex_width-1:i*vertex_width], getVertex_60[(i+1)*vertex_width-1:i*vertex_width], getVertex_61[(i+1)*vertex_width-1:i*vertex_width], getVertex_62[(i+1)*vertex_width-1:i*vertex_width], getVertex_63[(i+1)*vertex_width-1:i*vertex_width]} = data_in[(folding_factor-i)*vertex_width*64-1:(folding_factor-i-1)*vertex_width*64];
   end
endgenerate
	
//assign data_o = {vertex_0[3:0], vertex_1[3:0], vertex_2[3:0], vertex_3[3:0], vertex_4[3:0], vertex_5[3:0], vertex_6[3:0], vertex_7[3:0], vertex_8[3:0], vertex_9[3:0], vertex_10[3:0], vertex_11[3:0], vertex_12[3:0], vertex_13[3:0], vertex_14[3:0], vertex_15[3:0], vertex_16[3:0], vertex_17[3:0], vertex_18[3:0], vertex_19[3:0], vertex_20[3:0], vertex_21[3:0], vertex_22[3:0], vertex_23[3:0], vertex_24[3:0], vertex_25[3:0], vertex_26[3:0], vertex_27[3:0], vertex_28[3:0], vertex_29[3:0], vertex_30[3:0], vertex_31[3:0], vertex_32[3:0], vertex_33[3:0], vertex_34[3:0], vertex_35[3:0], vertex_36[3:0], vertex_37[3:0], vertex_38[3:0], vertex_39[3:0], vertex_40[3:0], vertex_41[3:0], vertex_42[3:0], vertex_43[3:0], vertex_44[3:0], vertex_45[3:0], vertex_46[3:0], vertex_47[3:0], vertex_48[3:0], vertex_49[3:0], vertex_50[3:0], vertex_51[3:0], vertex_52[3:0], vertex_53[3:0], vertex_54[3:0], vertex_55[3:0], vertex_56[3:0], vertex_57[3:0], vertex_58[3:0], vertex_59[3:0], vertex_60[3:0], vertex_61[3:0], vertex_62[3:0], vertex_63[3:0], vertex_0[7:4], vertex_1[7:4], vertex_2[7:4], vertex_3[7:4], vertex_4[7:4], vertex_5[7:4], vertex_6[7:4], vertex_7[7:4], vertex_8[7:4], vertex_9[7:4], vertex_10[7:4], vertex_11[7:4], vertex_12[7:4], vertex_13[7:4], vertex_14[7:4], vertex_15[7:4], vertex_16[7:4], vertex_17[7:4], vertex_18[7:4], vertex_19[7:4], vertex_20[7:4], vertex_21[7:4], vertex_22[7:4], vertex_23[7:4], vertex_24[7:4], vertex_25[7:4], vertex_26[7:4], vertex_27[7:4], vertex_28[7:4], vertex_29[7:4], vertex_30[7:4], vertex_31[7:4], vertex_32[7:4], vertex_33[7:4], vertex_34[7:4], vertex_35[7:4], vertex_36[7:4], vertex_37[7:4], vertex_38[7:4], vertex_39[7:4], vertex_40[7:4], vertex_41[7:4], vertex_42[7:4], vertex_43[7:4], vertex_44[7:4], vertex_45[7:4], vertex_46[7:4], vertex_47[7:4], vertex_48[7:4], vertex_49[7:4], vertex_50[7:4], vertex_51[7:4], vertex_52[7:4], vertex_53[7:4], vertex_54[7:4], vertex_55[7:4], vertex_56[7:4], vertex_57[7:4], vertex_58[7:4], vertex_59[7:4], vertex_60[7:4], vertex_61[7:4], vertex_62[7:4], vertex_63[7:4], vertex_0[11:8], vertex_1[11:8], vertex_2[11:8], vertex_3[11:8], vertex_4[11:8], vertex_5[11:8], vertex_6[11:8], vertex_7[11:8], vertex_8[11:8], vertex_9[11:8], vertex_10[11:8], vertex_11[11:8], vertex_12[11:8], vertex_13[11:8], vertex_14[11:8], vertex_15[11:8], vertex_16[11:8], vertex_17[11:8], vertex_18[11:8], vertex_19[11:8], vertex_20[11:8], vertex_21[11:8], vertex_22[11:8], vertex_23[11:8], vertex_24[11:8], vertex_25[11:8], vertex_26[11:8], vertex_27[11:8], vertex_28[11:8], vertex_29[11:8], vertex_30[11:8], vertex_31[11:8], vertex_32[11:8], vertex_33[11:8], vertex_34[11:8], vertex_35[11:8], vertex_36[11:8], vertex_37[11:8], vertex_38[11:8], vertex_39[11:8], vertex_40[11:8], vertex_41[11:8], vertex_42[11:8], vertex_43[11:8], vertex_44[11:8], vertex_45[11:8], vertex_46[11:8], vertex_47[11:8], vertex_48[11:8], vertex_49[11:8], vertex_50[11:8], vertex_51[11:8], vertex_52[11:8], vertex_53[11:8], vertex_54[11:8], vertex_55[11:8], vertex_56[11:8], vertex_57[11:8], vertex_58[11:8], vertex_59[11:8], vertex_60[11:8], vertex_61[11:8], vertex_62[11:8], vertex_63[11:8], vertex_0[15:12], vertex_1[15:12], vertex_2[15:12], vertex_3[15:12], vertex_4[15:12], vertex_5[15:12], vertex_6[15:12], vertex_7[15:12], vertex_8[15:12], vertex_9[15:12], vertex_10[15:12], vertex_11[15:12], vertex_12[15:12], vertex_13[15:12], vertex_14[15:12], vertex_15[15:12], vertex_16[15:12], vertex_17[15:12], vertex_18[15:12], vertex_19[15:12], vertex_20[15:12], vertex_21[15:12], vertex_22[15:12], vertex_23[15:12], vertex_24[15:12], vertex_25[15:12], vertex_26[15:12], vertex_27[15:12], vertex_28[15:12], vertex_29[15:12], vertex_30[15:12], vertex_31[15:12], vertex_32[15:12], vertex_33[15:12], vertex_34[15:12], vertex_35[15:12], vertex_36[15:12], vertex_37[15:12], vertex_38[15:12], vertex_39[15:12], vertex_40[15:12], vertex_41[15:12], vertex_42[15:12], vertex_43[15:12], vertex_44[15:12], vertex_45[15:12], vertex_46[15:12], vertex_47[15:12], vertex_48[15:12], vertex_49[15:12], vertex_50[15:12], vertex_51[15:12], vertex_52[15:12], vertex_53[15:12], vertex_54[15:12], vertex_55[15:12], vertex_56[15:12], vertex_57[15:12], vertex_58[15:12], vertex_59[15:12], vertex_60[15:12], vertex_61[15:12], vertex_62[15:12], vertex_63[15:12]};

//assign {getVertex_0[3:0], getVertex_1[3:0], getVertex_2[3:0], getVertex_3[3:0], getVertex_4[3:0], getVertex_5[3:0], getVertex_6[3:0], getVertex_7[3:0], getVertex_8[3:0], getVertex_9[3:0], getVertex_10[3:0], getVertex_11[3:0], getVertex_12[3:0], getVertex_13[3:0], getVertex_14[3:0], getVertex_15[3:0], getVertex_16[3:0], getVertex_17[3:0], getVertex_18[3:0], getVertex_19[3:0], getVertex_20[3:0], getVertex_21[3:0], getVertex_22[3:0], getVertex_23[3:0], getVertex_24[3:0], getVertex_25[3:0], getVertex_26[3:0], getVertex_27[3:0], getVertex_28[3:0], getVertex_29[3:0], getVertex_30[3:0], getVertex_31[3:0], getVertex_32[3:0], getVertex_33[3:0], getVertex_34[3:0], getVertex_35[3:0], getVertex_36[3:0], getVertex_37[3:0], getVertex_38[3:0], getVertex_39[3:0], getVertex_40[3:0], getVertex_41[3:0], getVertex_42[3:0], getVertex_43[3:0], getVertex_44[3:0], getVertex_45[3:0], getVertex_46[3:0], getVertex_47[3:0], getVertex_48[3:0], getVertex_49[3:0], getVertex_50[3:0], getVertex_51[3:0], getVertex_52[3:0], getVertex_53[3:0], getVertex_54[3:0], getVertex_55[3:0], getVertex_56[3:0], getVertex_57[3:0], getVertex_58[3:0], getVertex_59[3:0], getVertex_60[3:0], getVertex_61[3:0], getVertex_62[3:0], getVertex_63[3:0], getVertex_0[7:4], getVertex_1[7:4], getVertex_2[7:4], getVertex_3[7:4], getVertex_4[7:4], getVertex_5[7:4], getVertex_6[7:4], getVertex_7[7:4], getVertex_8[7:4], getVertex_9[7:4], getVertex_10[7:4], getVertex_11[7:4], getVertex_12[7:4], getVertex_13[7:4], getVertex_14[7:4], getVertex_15[7:4], getVertex_16[7:4], getVertex_17[7:4], getVertex_18[7:4], getVertex_19[7:4], getVertex_20[7:4], getVertex_21[7:4], getVertex_22[7:4], getVertex_23[7:4], getVertex_24[7:4], getVertex_25[7:4], getVertex_26[7:4], getVertex_27[7:4], getVertex_28[7:4], getVertex_29[7:4], getVertex_30[7:4], getVertex_31[7:4], getVertex_32[7:4], getVertex_33[7:4], getVertex_34[7:4], getVertex_35[7:4], getVertex_36[7:4], getVertex_37[7:4], getVertex_38[7:4], getVertex_39[7:4], getVertex_40[7:4], getVertex_41[7:4], getVertex_42[7:4], getVertex_43[7:4], getVertex_44[7:4], getVertex_45[7:4], getVertex_46[7:4], getVertex_47[7:4], getVertex_48[7:4], getVertex_49[7:4], getVertex_50[7:4], getVertex_51[7:4], getVertex_52[7:4], getVertex_53[7:4], getVertex_54[7:4], getVertex_55[7:4], getVertex_56[7:4], getVertex_57[7:4], getVertex_58[7:4], getVertex_59[7:4], getVertex_60[7:4], getVertex_61[7:4], getVertex_62[7:4], getVertex_63[7:4], getVertex_0[11:8], getVertex_1[11:8], getVertex_2[11:8], getVertex_3[11:8], getVertex_4[11:8], getVertex_5[11:8], getVertex_6[11:8], getVertex_7[11:8], getVertex_8[11:8], getVertex_9[11:8], getVertex_10[11:8], getVertex_11[11:8], getVertex_12[11:8], getVertex_13[11:8], getVertex_14[11:8], getVertex_15[11:8], getVertex_16[11:8], getVertex_17[11:8], getVertex_18[11:8], getVertex_19[11:8], getVertex_20[11:8], getVertex_21[11:8], getVertex_22[11:8], getVertex_23[11:8], getVertex_24[11:8], getVertex_25[11:8], getVertex_26[11:8], getVertex_27[11:8], getVertex_28[11:8], getVertex_29[11:8], getVertex_30[11:8], getVertex_31[11:8], getVertex_32[11:8], getVertex_33[11:8], getVertex_34[11:8], getVertex_35[11:8], getVertex_36[11:8], getVertex_37[11:8], getVertex_38[11:8], getVertex_39[11:8], getVertex_40[11:8], getVertex_41[11:8], getVertex_42[11:8], getVertex_43[11:8], getVertex_44[11:8], getVertex_45[11:8], getVertex_46[11:8], getVertex_47[11:8], getVertex_48[11:8], getVertex_49[11:8], getVertex_50[11:8], getVertex_51[11:8], getVertex_52[11:8], getVertex_53[11:8], getVertex_54[11:8], getVertex_55[11:8], getVertex_56[11:8], getVertex_57[11:8], getVertex_58[11:8], getVertex_59[11:8], getVertex_60[11:8], getVertex_61[11:8], getVertex_62[11:8], getVertex_63[11:8], getVertex_0[15:12], getVertex_1[15:12], getVertex_2[15:12], getVertex_3[15:12], getVertex_4[15:12], getVertex_5[15:12], getVertex_6[15:12], getVertex_7[15:12], getVertex_8[15:12], getVertex_9[15:12], getVertex_10[15:12], getVertex_11[15:12], getVertex_12[15:12], getVertex_13[15:12], getVertex_14[15:12], getVertex_15[15:12], getVertex_16[15:12], getVertex_17[15:12], getVertex_18[15:12], getVertex_19[15:12], getVertex_20[15:12], getVertex_21[15:12], getVertex_22[15:12], getVertex_23[15:12], getVertex_24[15:12], getVertex_25[15:12], getVertex_26[15:12], getVertex_27[15:12], getVertex_28[15:12], getVertex_29[15:12], getVertex_30[15:12], getVertex_31[15:12], getVertex_32[15:12], getVertex_33[15:12], getVertex_34[15:12], getVertex_35[15:12], getVertex_36[15:12], getVertex_37[15:12], getVertex_38[15:12], getVertex_39[15:12], getVertex_40[15:12], getVertex_41[15:12], getVertex_42[15:12], getVertex_43[15:12], getVertex_44[15:12], getVertex_45[15:12], getVertex_46[15:12], getVertex_47[15:12], getVertex_48[15:12], getVertex_49[15:12], getVertex_50[15:12], getVertex_51[15:12], getVertex_52[15:12], getVertex_53[15:12], getVertex_54[15:12], getVertex_55[15:12], getVertex_56[15:12], getVertex_57[15:12], getVertex_58[15:12], getVertex_59[15:12], getVertex_60[15:12], getVertex_61[15:12], getVertex_62[15:12], getVertex_63[15:12]} = data_in;


myNetworkYatish Net
			(
			.CLK(clk)
			,.RST_N(rst_n)
			, .send_ports_0_putFlit_flit_in(send_ports_0_putFlit_flit_in)
			, .EN_send_ports_0_putFlit(EN_send_ports_0_putFlit)
			, .EN_send_ports_0_getNonFullVCs(1'b1)
			, .send_ports_0_getNonFullVCs(send_ports_0_getNonFullVCs)
			, .recv_ports_0_getFlit(recv_ports_0_getFlit)
			, .EN_recv_ports_0_getFlit(EN_recv_ports_0_getFlit)
			, .EN_recv_ports_0_putNonFullVCs(1'b1)
			, .recv_ports_0_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_0_getRecvPortID(recv_ports_info_0_getRecvPortID)
			

			, .send_ports_1_putFlit_flit_in(send_ports_1_putFlit_flit_in)
			, .EN_send_ports_1_putFlit(EN_send_ports_1_putFlit)
			, .EN_send_ports_1_getNonFullVCs(1'b1)
			, .send_ports_1_getNonFullVCs(send_ports_1_getNonFullVCs)
			, .recv_ports_1_getFlit(recv_ports_1_getFlit)
			, .EN_recv_ports_1_getFlit(EN_recv_ports_1_getFlit)
			, .EN_recv_ports_1_putNonFullVCs(1'b1)
			, .recv_ports_1_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_1_getRecvPortID(recv_ports_info_1_getRecvPortID)
			

			, .send_ports_2_putFlit_flit_in(send_ports_2_putFlit_flit_in)
			, .EN_send_ports_2_putFlit(EN_send_ports_2_putFlit)
			, .EN_send_ports_2_getNonFullVCs(1'b1)
			, .send_ports_2_getNonFullVCs(send_ports_2_getNonFullVCs)
			, .recv_ports_2_getFlit(recv_ports_2_getFlit)
			, .EN_recv_ports_2_getFlit(EN_recv_ports_2_getFlit)
			, .EN_recv_ports_2_putNonFullVCs(1'b1)
			, .recv_ports_2_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_2_getRecvPortID(recv_ports_info_2_getRecvPortID)
			

			, .send_ports_3_putFlit_flit_in(send_ports_3_putFlit_flit_in)
			, .EN_send_ports_3_putFlit(EN_send_ports_3_putFlit)
			, .EN_send_ports_3_getNonFullVCs(1'b1)
			, .send_ports_3_getNonFullVCs(send_ports_3_getNonFullVCs)
			, .recv_ports_3_getFlit(recv_ports_3_getFlit)
			, .EN_recv_ports_3_getFlit(EN_recv_ports_3_getFlit)
			, .EN_recv_ports_3_putNonFullVCs(1'b1)
			, .recv_ports_3_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_3_getRecvPortID(recv_ports_info_3_getRecvPortID)
			

			, .send_ports_4_putFlit_flit_in(send_ports_4_putFlit_flit_in)
			, .EN_send_ports_4_putFlit(EN_send_ports_4_putFlit)
			, .EN_send_ports_4_getNonFullVCs(1'b1)
			, .send_ports_4_getNonFullVCs(send_ports_4_getNonFullVCs)
			, .recv_ports_4_getFlit(recv_ports_4_getFlit)
			, .EN_recv_ports_4_getFlit(EN_recv_ports_4_getFlit)
			, .EN_recv_ports_4_putNonFullVCs(1'b1)
			, .recv_ports_4_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_4_getRecvPortID(recv_ports_info_4_getRecvPortID)
			

			, .send_ports_5_putFlit_flit_in(send_ports_5_putFlit_flit_in)
			, .EN_send_ports_5_putFlit(EN_send_ports_5_putFlit)
			, .EN_send_ports_5_getNonFullVCs(1'b1)
			, .send_ports_5_getNonFullVCs(send_ports_5_getNonFullVCs)
			, .recv_ports_5_getFlit(recv_ports_5_getFlit)
			, .EN_recv_ports_5_getFlit(EN_recv_ports_5_getFlit)
			, .EN_recv_ports_5_putNonFullVCs(1'b1)
			, .recv_ports_5_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_5_getRecvPortID(recv_ports_info_5_getRecvPortID)
			

			, .send_ports_6_putFlit_flit_in(send_ports_6_putFlit_flit_in)
			, .EN_send_ports_6_putFlit(EN_send_ports_6_putFlit)
			, .EN_send_ports_6_getNonFullVCs(1'b1)
			, .send_ports_6_getNonFullVCs(send_ports_6_getNonFullVCs)
			, .recv_ports_6_getFlit(recv_ports_6_getFlit)
			, .EN_recv_ports_6_getFlit(EN_recv_ports_6_getFlit)
			, .EN_recv_ports_6_putNonFullVCs(1'b1)
			, .recv_ports_6_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_6_getRecvPortID(recv_ports_info_6_getRecvPortID)
			

			, .send_ports_7_putFlit_flit_in(send_ports_7_putFlit_flit_in)
			, .EN_send_ports_7_putFlit(EN_send_ports_7_putFlit)
			, .EN_send_ports_7_getNonFullVCs(1'b1)
			, .send_ports_7_getNonFullVCs(send_ports_7_getNonFullVCs)
			, .recv_ports_7_getFlit(recv_ports_7_getFlit)
			, .EN_recv_ports_7_getFlit(EN_recv_ports_7_getFlit)
			, .EN_recv_ports_7_putNonFullVCs(1'b1)
			, .recv_ports_7_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_7_getRecvPortID(recv_ports_info_7_getRecvPortID)
			

			, .send_ports_8_putFlit_flit_in(send_ports_8_putFlit_flit_in)
			, .EN_send_ports_8_putFlit(EN_send_ports_8_putFlit)
			, .EN_send_ports_8_getNonFullVCs(1'b1)
			, .send_ports_8_getNonFullVCs(send_ports_8_getNonFullVCs)
			, .recv_ports_8_getFlit(recv_ports_8_getFlit)
			, .EN_recv_ports_8_getFlit(EN_recv_ports_8_getFlit)
			, .EN_recv_ports_8_putNonFullVCs(1'b1)
			, .recv_ports_8_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_8_getRecvPortID(recv_ports_info_8_getRecvPortID)
			

			, .send_ports_9_putFlit_flit_in(send_ports_9_putFlit_flit_in)
			, .EN_send_ports_9_putFlit(EN_send_ports_9_putFlit)
			, .EN_send_ports_9_getNonFullVCs(1'b1)
			, .send_ports_9_getNonFullVCs(send_ports_9_getNonFullVCs)
			, .recv_ports_9_getFlit(recv_ports_9_getFlit)
			, .EN_recv_ports_9_getFlit(EN_recv_ports_9_getFlit)
			, .EN_recv_ports_9_putNonFullVCs(1'b1)
			, .recv_ports_9_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_9_getRecvPortID(recv_ports_info_9_getRecvPortID)
			

			, .send_ports_10_putFlit_flit_in(send_ports_10_putFlit_flit_in)
			, .EN_send_ports_10_putFlit(EN_send_ports_10_putFlit)
			, .EN_send_ports_10_getNonFullVCs(1'b1)
			, .send_ports_10_getNonFullVCs(send_ports_10_getNonFullVCs)
			, .recv_ports_10_getFlit(recv_ports_10_getFlit)
			, .EN_recv_ports_10_getFlit(EN_recv_ports_10_getFlit)
			, .EN_recv_ports_10_putNonFullVCs(1'b1)
			, .recv_ports_10_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_10_getRecvPortID(recv_ports_info_10_getRecvPortID)
			

			, .send_ports_11_putFlit_flit_in(send_ports_11_putFlit_flit_in)
			, .EN_send_ports_11_putFlit(EN_send_ports_11_putFlit)
			, .EN_send_ports_11_getNonFullVCs(1'b1)
			, .send_ports_11_getNonFullVCs(send_ports_11_getNonFullVCs)
			, .recv_ports_11_getFlit(recv_ports_11_getFlit)
			, .EN_recv_ports_11_getFlit(EN_recv_ports_11_getFlit)
			, .EN_recv_ports_11_putNonFullVCs(1'b1)
			, .recv_ports_11_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_11_getRecvPortID(recv_ports_info_11_getRecvPortID)
			

			, .send_ports_12_putFlit_flit_in(send_ports_12_putFlit_flit_in)
			, .EN_send_ports_12_putFlit(EN_send_ports_12_putFlit)
			, .EN_send_ports_12_getNonFullVCs(1'b1)
			, .send_ports_12_getNonFullVCs(send_ports_12_getNonFullVCs)
			, .recv_ports_12_getFlit(recv_ports_12_getFlit)
			, .EN_recv_ports_12_getFlit(EN_recv_ports_12_getFlit)
			, .EN_recv_ports_12_putNonFullVCs(1'b1)
			, .recv_ports_12_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_12_getRecvPortID(recv_ports_info_12_getRecvPortID)
			

			, .send_ports_13_putFlit_flit_in(send_ports_13_putFlit_flit_in)
			, .EN_send_ports_13_putFlit(EN_send_ports_13_putFlit)
			, .EN_send_ports_13_getNonFullVCs(1'b1)
			, .send_ports_13_getNonFullVCs(send_ports_13_getNonFullVCs)
			, .recv_ports_13_getFlit(recv_ports_13_getFlit)
			, .EN_recv_ports_13_getFlit(EN_recv_ports_13_getFlit)
			, .EN_recv_ports_13_putNonFullVCs(1'b1)
			, .recv_ports_13_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_13_getRecvPortID(recv_ports_info_13_getRecvPortID)
			

			, .send_ports_14_putFlit_flit_in(send_ports_14_putFlit_flit_in)
			, .EN_send_ports_14_putFlit(EN_send_ports_14_putFlit)
			, .EN_send_ports_14_getNonFullVCs(1'b1)
			, .send_ports_14_getNonFullVCs(send_ports_14_getNonFullVCs)
			, .recv_ports_14_getFlit(recv_ports_14_getFlit)
			, .EN_recv_ports_14_getFlit(EN_recv_ports_14_getFlit)
			, .EN_recv_ports_14_putNonFullVCs(1'b1)
			, .recv_ports_14_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_14_getRecvPortID(recv_ports_info_14_getRecvPortID)
			

			, .send_ports_15_putFlit_flit_in(send_ports_15_putFlit_flit_in)
			, .EN_send_ports_15_putFlit(EN_send_ports_15_putFlit)
			, .EN_send_ports_15_getNonFullVCs(1'b1)
			, .send_ports_15_getNonFullVCs(send_ports_15_getNonFullVCs)
			, .recv_ports_15_getFlit(recv_ports_15_getFlit)
			, .EN_recv_ports_15_getFlit(EN_recv_ports_15_getFlit)
			, .EN_recv_ports_15_putNonFullVCs(1'b1)
			, .recv_ports_15_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_15_getRecvPortID(recv_ports_info_15_getRecvPortID)
			

			, .send_ports_16_putFlit_flit_in(send_ports_16_putFlit_flit_in)
			, .EN_send_ports_16_putFlit(EN_send_ports_16_putFlit)
			, .EN_send_ports_16_getNonFullVCs(1'b1)
			, .send_ports_16_getNonFullVCs(send_ports_16_getNonFullVCs)
			, .recv_ports_16_getFlit(recv_ports_16_getFlit)
			, .EN_recv_ports_16_getFlit(EN_recv_ports_16_getFlit)
			, .EN_recv_ports_16_putNonFullVCs(1'b1)
			, .recv_ports_16_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_16_getRecvPortID(recv_ports_info_16_getRecvPortID)
			

			, .send_ports_17_putFlit_flit_in(send_ports_17_putFlit_flit_in)
			, .EN_send_ports_17_putFlit(EN_send_ports_17_putFlit)
			, .EN_send_ports_17_getNonFullVCs(1'b1)
			, .send_ports_17_getNonFullVCs(send_ports_17_getNonFullVCs)
			, .recv_ports_17_getFlit(recv_ports_17_getFlit)
			, .EN_recv_ports_17_getFlit(EN_recv_ports_17_getFlit)
			, .EN_recv_ports_17_putNonFullVCs(1'b1)
			, .recv_ports_17_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_17_getRecvPortID(recv_ports_info_17_getRecvPortID)
			

			, .send_ports_18_putFlit_flit_in(send_ports_18_putFlit_flit_in)
			, .EN_send_ports_18_putFlit(EN_send_ports_18_putFlit)
			, .EN_send_ports_18_getNonFullVCs(1'b1)
			, .send_ports_18_getNonFullVCs(send_ports_18_getNonFullVCs)
			, .recv_ports_18_getFlit(recv_ports_18_getFlit)
			, .EN_recv_ports_18_getFlit(EN_recv_ports_18_getFlit)
			, .EN_recv_ports_18_putNonFullVCs(1'b1)
			, .recv_ports_18_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_18_getRecvPortID(recv_ports_info_18_getRecvPortID)
			

			, .send_ports_19_putFlit_flit_in(send_ports_19_putFlit_flit_in)
			, .EN_send_ports_19_putFlit(EN_send_ports_19_putFlit)
			, .EN_send_ports_19_getNonFullVCs(1'b1)
			, .send_ports_19_getNonFullVCs(send_ports_19_getNonFullVCs)
			, .recv_ports_19_getFlit(recv_ports_19_getFlit)
			, .EN_recv_ports_19_getFlit(EN_recv_ports_19_getFlit)
			, .EN_recv_ports_19_putNonFullVCs(1'b1)
			, .recv_ports_19_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_19_getRecvPortID(recv_ports_info_19_getRecvPortID)
			

			, .send_ports_20_putFlit_flit_in(send_ports_20_putFlit_flit_in)
			, .EN_send_ports_20_putFlit(EN_send_ports_20_putFlit)
			, .EN_send_ports_20_getNonFullVCs(1'b1)
			, .send_ports_20_getNonFullVCs(send_ports_20_getNonFullVCs)
			, .recv_ports_20_getFlit(recv_ports_20_getFlit)
			, .EN_recv_ports_20_getFlit(EN_recv_ports_20_getFlit)
			, .EN_recv_ports_20_putNonFullVCs(1'b1)
			, .recv_ports_20_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_20_getRecvPortID(recv_ports_info_20_getRecvPortID)
			

			, .send_ports_21_putFlit_flit_in(send_ports_21_putFlit_flit_in)
			, .EN_send_ports_21_putFlit(EN_send_ports_21_putFlit)
			, .EN_send_ports_21_getNonFullVCs(1'b1)
			, .send_ports_21_getNonFullVCs(send_ports_21_getNonFullVCs)
			, .recv_ports_21_getFlit(recv_ports_21_getFlit)
			, .EN_recv_ports_21_getFlit(EN_recv_ports_21_getFlit)
			, .EN_recv_ports_21_putNonFullVCs(1'b1)
			, .recv_ports_21_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_21_getRecvPortID(recv_ports_info_21_getRecvPortID)
			

			, .send_ports_22_putFlit_flit_in(send_ports_22_putFlit_flit_in)
			, .EN_send_ports_22_putFlit(EN_send_ports_22_putFlit)
			, .EN_send_ports_22_getNonFullVCs(1'b1)
			, .send_ports_22_getNonFullVCs(send_ports_22_getNonFullVCs)
			, .recv_ports_22_getFlit(recv_ports_22_getFlit)
			, .EN_recv_ports_22_getFlit(EN_recv_ports_22_getFlit)
			, .EN_recv_ports_22_putNonFullVCs(1'b1)
			, .recv_ports_22_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_22_getRecvPortID(recv_ports_info_22_getRecvPortID)
			

			, .send_ports_23_putFlit_flit_in(send_ports_23_putFlit_flit_in)
			, .EN_send_ports_23_putFlit(EN_send_ports_23_putFlit)
			, .EN_send_ports_23_getNonFullVCs(1'b1)
			, .send_ports_23_getNonFullVCs(send_ports_23_getNonFullVCs)
			, .recv_ports_23_getFlit(recv_ports_23_getFlit)
			, .EN_recv_ports_23_getFlit(EN_recv_ports_23_getFlit)
			, .EN_recv_ports_23_putNonFullVCs(1'b1)
			, .recv_ports_23_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_23_getRecvPortID(recv_ports_info_23_getRecvPortID)
			

			, .send_ports_24_putFlit_flit_in(send_ports_24_putFlit_flit_in)
			, .EN_send_ports_24_putFlit(EN_send_ports_24_putFlit)
			, .EN_send_ports_24_getNonFullVCs(1'b1)
			, .send_ports_24_getNonFullVCs(send_ports_24_getNonFullVCs)
			, .recv_ports_24_getFlit(recv_ports_24_getFlit)
			, .EN_recv_ports_24_getFlit(EN_recv_ports_24_getFlit)
			, .EN_recv_ports_24_putNonFullVCs(1'b1)
			, .recv_ports_24_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_24_getRecvPortID(recv_ports_info_24_getRecvPortID)
			

			, .send_ports_25_putFlit_flit_in(send_ports_25_putFlit_flit_in)
			, .EN_send_ports_25_putFlit(EN_send_ports_25_putFlit)
			, .EN_send_ports_25_getNonFullVCs(1'b1)
			, .send_ports_25_getNonFullVCs(send_ports_25_getNonFullVCs)
			, .recv_ports_25_getFlit(recv_ports_25_getFlit)
			, .EN_recv_ports_25_getFlit(EN_recv_ports_25_getFlit)
			, .EN_recv_ports_25_putNonFullVCs(1'b1)
			, .recv_ports_25_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_25_getRecvPortID(recv_ports_info_25_getRecvPortID)
			

			, .send_ports_26_putFlit_flit_in(send_ports_26_putFlit_flit_in)
			, .EN_send_ports_26_putFlit(EN_send_ports_26_putFlit)
			, .EN_send_ports_26_getNonFullVCs(1'b1)
			, .send_ports_26_getNonFullVCs(send_ports_26_getNonFullVCs)
			, .recv_ports_26_getFlit(recv_ports_26_getFlit)
			, .EN_recv_ports_26_getFlit(EN_recv_ports_26_getFlit)
			, .EN_recv_ports_26_putNonFullVCs(1'b1)
			, .recv_ports_26_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_26_getRecvPortID(recv_ports_info_26_getRecvPortID)
			

			, .send_ports_27_putFlit_flit_in(send_ports_27_putFlit_flit_in)
			, .EN_send_ports_27_putFlit(EN_send_ports_27_putFlit)
			, .EN_send_ports_27_getNonFullVCs(1'b1)
			, .send_ports_27_getNonFullVCs(send_ports_27_getNonFullVCs)
			, .recv_ports_27_getFlit(recv_ports_27_getFlit)
			, .EN_recv_ports_27_getFlit(EN_recv_ports_27_getFlit)
			, .EN_recv_ports_27_putNonFullVCs(1'b1)
			, .recv_ports_27_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_27_getRecvPortID(recv_ports_info_27_getRecvPortID)
			

			, .send_ports_28_putFlit_flit_in(send_ports_28_putFlit_flit_in)
			, .EN_send_ports_28_putFlit(EN_send_ports_28_putFlit)
			, .EN_send_ports_28_getNonFullVCs(1'b1)
			, .send_ports_28_getNonFullVCs(send_ports_28_getNonFullVCs)
			, .recv_ports_28_getFlit(recv_ports_28_getFlit)
			, .EN_recv_ports_28_getFlit(EN_recv_ports_28_getFlit)
			, .EN_recv_ports_28_putNonFullVCs(1'b1)
			, .recv_ports_28_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_28_getRecvPortID(recv_ports_info_28_getRecvPortID)
			

			, .send_ports_29_putFlit_flit_in(send_ports_29_putFlit_flit_in)
			, .EN_send_ports_29_putFlit(EN_send_ports_29_putFlit)
			, .EN_send_ports_29_getNonFullVCs(1'b1)
			, .send_ports_29_getNonFullVCs(send_ports_29_getNonFullVCs)
			, .recv_ports_29_getFlit(recv_ports_29_getFlit)
			, .EN_recv_ports_29_getFlit(EN_recv_ports_29_getFlit)
			, .EN_recv_ports_29_putNonFullVCs(1'b1)
			, .recv_ports_29_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_29_getRecvPortID(recv_ports_info_29_getRecvPortID)
			

			, .send_ports_30_putFlit_flit_in(send_ports_30_putFlit_flit_in)
			, .EN_send_ports_30_putFlit(EN_send_ports_30_putFlit)
			, .EN_send_ports_30_getNonFullVCs(1'b1)
			, .send_ports_30_getNonFullVCs(send_ports_30_getNonFullVCs)
			, .recv_ports_30_getFlit(recv_ports_30_getFlit)
			, .EN_recv_ports_30_getFlit(EN_recv_ports_30_getFlit)
			, .EN_recv_ports_30_putNonFullVCs(1'b1)
			, .recv_ports_30_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_30_getRecvPortID(recv_ports_info_30_getRecvPortID)
			

			, .send_ports_31_putFlit_flit_in(send_ports_31_putFlit_flit_in)
			, .EN_send_ports_31_putFlit(EN_send_ports_31_putFlit)
			, .EN_send_ports_31_getNonFullVCs(1'b1)
			, .send_ports_31_getNonFullVCs(send_ports_31_getNonFullVCs)
			, .recv_ports_31_getFlit(recv_ports_31_getFlit)
			, .EN_recv_ports_31_getFlit(EN_recv_ports_31_getFlit)
			, .EN_recv_ports_31_putNonFullVCs(1'b1)
			, .recv_ports_31_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_31_getRecvPortID(recv_ports_info_31_getRecvPortID)
			

			, .send_ports_32_putFlit_flit_in(send_ports_32_putFlit_flit_in)
			, .EN_send_ports_32_putFlit(EN_send_ports_32_putFlit)
			, .EN_send_ports_32_getNonFullVCs(1'b1)
			, .send_ports_32_getNonFullVCs(send_ports_32_getNonFullVCs)
			, .recv_ports_32_getFlit(recv_ports_32_getFlit)
			, .EN_recv_ports_32_getFlit(EN_recv_ports_32_getFlit)
			, .EN_recv_ports_32_putNonFullVCs(1'b1)
			, .recv_ports_32_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_32_getRecvPortID(recv_ports_info_32_getRecvPortID)
			

			, .send_ports_33_putFlit_flit_in(send_ports_33_putFlit_flit_in)
			, .EN_send_ports_33_putFlit(EN_send_ports_33_putFlit)
			, .EN_send_ports_33_getNonFullVCs(1'b1)
			, .send_ports_33_getNonFullVCs(send_ports_33_getNonFullVCs)
			, .recv_ports_33_getFlit(recv_ports_33_getFlit)
			, .EN_recv_ports_33_getFlit(EN_recv_ports_33_getFlit)
			, .EN_recv_ports_33_putNonFullVCs(1'b1)
			, .recv_ports_33_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_33_getRecvPortID(recv_ports_info_33_getRecvPortID)
			

			, .send_ports_34_putFlit_flit_in(send_ports_34_putFlit_flit_in)
			, .EN_send_ports_34_putFlit(EN_send_ports_34_putFlit)
			, .EN_send_ports_34_getNonFullVCs(1'b1)
			, .send_ports_34_getNonFullVCs(send_ports_34_getNonFullVCs)
			, .recv_ports_34_getFlit(recv_ports_34_getFlit)
			, .EN_recv_ports_34_getFlit(EN_recv_ports_34_getFlit)
			, .EN_recv_ports_34_putNonFullVCs(1'b1)
			, .recv_ports_34_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_34_getRecvPortID(recv_ports_info_34_getRecvPortID)
			

			, .send_ports_35_putFlit_flit_in(send_ports_35_putFlit_flit_in)
			, .EN_send_ports_35_putFlit(EN_send_ports_35_putFlit)
			, .EN_send_ports_35_getNonFullVCs(1'b1)
			, .send_ports_35_getNonFullVCs(send_ports_35_getNonFullVCs)
			, .recv_ports_35_getFlit(recv_ports_35_getFlit)
			, .EN_recv_ports_35_getFlit(EN_recv_ports_35_getFlit)
			, .EN_recv_ports_35_putNonFullVCs(1'b1)
			, .recv_ports_35_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_35_getRecvPortID(recv_ports_info_35_getRecvPortID)
			

			, .send_ports_36_putFlit_flit_in(send_ports_36_putFlit_flit_in)
			, .EN_send_ports_36_putFlit(EN_send_ports_36_putFlit)
			, .EN_send_ports_36_getNonFullVCs(1'b1)
			, .send_ports_36_getNonFullVCs(send_ports_36_getNonFullVCs)
			, .recv_ports_36_getFlit(recv_ports_36_getFlit)
			, .EN_recv_ports_36_getFlit(EN_recv_ports_36_getFlit)
			, .EN_recv_ports_36_putNonFullVCs(1'b1)
			, .recv_ports_36_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_36_getRecvPortID(recv_ports_info_36_getRecvPortID)
			

			, .send_ports_37_putFlit_flit_in(send_ports_37_putFlit_flit_in)
			, .EN_send_ports_37_putFlit(EN_send_ports_37_putFlit)
			, .EN_send_ports_37_getNonFullVCs(1'b1)
			, .send_ports_37_getNonFullVCs(send_ports_37_getNonFullVCs)
			, .recv_ports_37_getFlit(recv_ports_37_getFlit)
			, .EN_recv_ports_37_getFlit(EN_recv_ports_37_getFlit)
			, .EN_recv_ports_37_putNonFullVCs(1'b1)
			, .recv_ports_37_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_37_getRecvPortID(recv_ports_info_37_getRecvPortID)
			

			, .send_ports_38_putFlit_flit_in(send_ports_38_putFlit_flit_in)
			, .EN_send_ports_38_putFlit(EN_send_ports_38_putFlit)
			, .EN_send_ports_38_getNonFullVCs(1'b1)
			, .send_ports_38_getNonFullVCs(send_ports_38_getNonFullVCs)
			, .recv_ports_38_getFlit(recv_ports_38_getFlit)
			, .EN_recv_ports_38_getFlit(EN_recv_ports_38_getFlit)
			, .EN_recv_ports_38_putNonFullVCs(1'b1)
			, .recv_ports_38_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_38_getRecvPortID(recv_ports_info_38_getRecvPortID)
			

			, .send_ports_39_putFlit_flit_in(send_ports_39_putFlit_flit_in)
			, .EN_send_ports_39_putFlit(EN_send_ports_39_putFlit)
			, .EN_send_ports_39_getNonFullVCs(1'b1)
			, .send_ports_39_getNonFullVCs(send_ports_39_getNonFullVCs)
			, .recv_ports_39_getFlit(recv_ports_39_getFlit)
			, .EN_recv_ports_39_getFlit(EN_recv_ports_39_getFlit)
			, .EN_recv_ports_39_putNonFullVCs(1'b1)
			, .recv_ports_39_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_39_getRecvPortID(recv_ports_info_39_getRecvPortID)
			

			, .send_ports_40_putFlit_flit_in(send_ports_40_putFlit_flit_in)
			, .EN_send_ports_40_putFlit(EN_send_ports_40_putFlit)
			, .EN_send_ports_40_getNonFullVCs(1'b1)
			, .send_ports_40_getNonFullVCs(send_ports_40_getNonFullVCs)
			, .recv_ports_40_getFlit(recv_ports_40_getFlit)
			, .EN_recv_ports_40_getFlit(EN_recv_ports_40_getFlit)
			, .EN_recv_ports_40_putNonFullVCs(1'b1)
			, .recv_ports_40_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_40_getRecvPortID(recv_ports_info_40_getRecvPortID)
			

			, .send_ports_41_putFlit_flit_in(send_ports_41_putFlit_flit_in)
			, .EN_send_ports_41_putFlit(EN_send_ports_41_putFlit)
			, .EN_send_ports_41_getNonFullVCs(1'b1)
			, .send_ports_41_getNonFullVCs(send_ports_41_getNonFullVCs)
			, .recv_ports_41_getFlit(recv_ports_41_getFlit)
			, .EN_recv_ports_41_getFlit(EN_recv_ports_41_getFlit)
			, .EN_recv_ports_41_putNonFullVCs(1'b1)
			, .recv_ports_41_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_41_getRecvPortID(recv_ports_info_41_getRecvPortID)
			

			, .send_ports_42_putFlit_flit_in(send_ports_42_putFlit_flit_in)
			, .EN_send_ports_42_putFlit(EN_send_ports_42_putFlit)
			, .EN_send_ports_42_getNonFullVCs(1'b1)
			, .send_ports_42_getNonFullVCs(send_ports_42_getNonFullVCs)
			, .recv_ports_42_getFlit(recv_ports_42_getFlit)
			, .EN_recv_ports_42_getFlit(EN_recv_ports_42_getFlit)
			, .EN_recv_ports_42_putNonFullVCs(1'b1)
			, .recv_ports_42_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_42_getRecvPortID(recv_ports_info_42_getRecvPortID)
			

			, .send_ports_43_putFlit_flit_in(send_ports_43_putFlit_flit_in)
			, .EN_send_ports_43_putFlit(EN_send_ports_43_putFlit)
			, .EN_send_ports_43_getNonFullVCs(1'b1)
			, .send_ports_43_getNonFullVCs(send_ports_43_getNonFullVCs)
			, .recv_ports_43_getFlit(recv_ports_43_getFlit)
			, .EN_recv_ports_43_getFlit(EN_recv_ports_43_getFlit)
			, .EN_recv_ports_43_putNonFullVCs(1'b1)
			, .recv_ports_43_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_43_getRecvPortID(recv_ports_info_43_getRecvPortID)
			

			, .send_ports_44_putFlit_flit_in(send_ports_44_putFlit_flit_in)
			, .EN_send_ports_44_putFlit(EN_send_ports_44_putFlit)
			, .EN_send_ports_44_getNonFullVCs(1'b1)
			, .send_ports_44_getNonFullVCs(send_ports_44_getNonFullVCs)
			, .recv_ports_44_getFlit(recv_ports_44_getFlit)
			, .EN_recv_ports_44_getFlit(EN_recv_ports_44_getFlit)
			, .EN_recv_ports_44_putNonFullVCs(1'b1)
			, .recv_ports_44_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_44_getRecvPortID(recv_ports_info_44_getRecvPortID)
			

			, .send_ports_45_putFlit_flit_in(send_ports_45_putFlit_flit_in)
			, .EN_send_ports_45_putFlit(EN_send_ports_45_putFlit)
			, .EN_send_ports_45_getNonFullVCs(1'b1)
			, .send_ports_45_getNonFullVCs(send_ports_45_getNonFullVCs)
			, .recv_ports_45_getFlit(recv_ports_45_getFlit)
			, .EN_recv_ports_45_getFlit(EN_recv_ports_45_getFlit)
			, .EN_recv_ports_45_putNonFullVCs(1'b1)
			, .recv_ports_45_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_45_getRecvPortID(recv_ports_info_45_getRecvPortID)
			

			, .send_ports_46_putFlit_flit_in(send_ports_46_putFlit_flit_in)
			, .EN_send_ports_46_putFlit(EN_send_ports_46_putFlit)
			, .EN_send_ports_46_getNonFullVCs(1'b1)
			, .send_ports_46_getNonFullVCs(send_ports_46_getNonFullVCs)
			, .recv_ports_46_getFlit(recv_ports_46_getFlit)
			, .EN_recv_ports_46_getFlit(EN_recv_ports_46_getFlit)
			, .EN_recv_ports_46_putNonFullVCs(1'b1)
			, .recv_ports_46_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_46_getRecvPortID(recv_ports_info_46_getRecvPortID)
			

			, .send_ports_47_putFlit_flit_in(send_ports_47_putFlit_flit_in)
			, .EN_send_ports_47_putFlit(EN_send_ports_47_putFlit)
			, .EN_send_ports_47_getNonFullVCs(1'b1)
			, .send_ports_47_getNonFullVCs(send_ports_47_getNonFullVCs)
			, .recv_ports_47_getFlit(recv_ports_47_getFlit)
			, .EN_recv_ports_47_getFlit(EN_recv_ports_47_getFlit)
			, .EN_recv_ports_47_putNonFullVCs(1'b1)
			, .recv_ports_47_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_47_getRecvPortID(recv_ports_info_47_getRecvPortID)
			

			, .send_ports_48_putFlit_flit_in(send_ports_48_putFlit_flit_in)
			, .EN_send_ports_48_putFlit(EN_send_ports_48_putFlit)
			, .EN_send_ports_48_getNonFullVCs(1'b1)
			, .send_ports_48_getNonFullVCs(send_ports_48_getNonFullVCs)
			, .recv_ports_48_getFlit(recv_ports_48_getFlit)
			, .EN_recv_ports_48_getFlit(EN_recv_ports_48_getFlit)
			, .EN_recv_ports_48_putNonFullVCs(1'b1)
			, .recv_ports_48_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_48_getRecvPortID(recv_ports_info_48_getRecvPortID)
			

			, .send_ports_49_putFlit_flit_in(send_ports_49_putFlit_flit_in)
			, .EN_send_ports_49_putFlit(EN_send_ports_49_putFlit)
			, .EN_send_ports_49_getNonFullVCs(1'b1)
			, .send_ports_49_getNonFullVCs(send_ports_49_getNonFullVCs)
			, .recv_ports_49_getFlit(recv_ports_49_getFlit)
			, .EN_recv_ports_49_getFlit(EN_recv_ports_49_getFlit)
			, .EN_recv_ports_49_putNonFullVCs(1'b1)
			, .recv_ports_49_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_49_getRecvPortID(recv_ports_info_49_getRecvPortID)
			

			, .send_ports_50_putFlit_flit_in(send_ports_50_putFlit_flit_in)
			, .EN_send_ports_50_putFlit(EN_send_ports_50_putFlit)
			, .EN_send_ports_50_getNonFullVCs(1'b1)
			, .send_ports_50_getNonFullVCs(send_ports_50_getNonFullVCs)
			, .recv_ports_50_getFlit(recv_ports_50_getFlit)
			, .EN_recv_ports_50_getFlit(EN_recv_ports_50_getFlit)
			, .EN_recv_ports_50_putNonFullVCs(1'b1)
			, .recv_ports_50_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_50_getRecvPortID(recv_ports_info_50_getRecvPortID)
			

			, .send_ports_51_putFlit_flit_in(send_ports_51_putFlit_flit_in)
			, .EN_send_ports_51_putFlit(EN_send_ports_51_putFlit)
			, .EN_send_ports_51_getNonFullVCs(1'b1)
			, .send_ports_51_getNonFullVCs(send_ports_51_getNonFullVCs)
			, .recv_ports_51_getFlit(recv_ports_51_getFlit)
			, .EN_recv_ports_51_getFlit(EN_recv_ports_51_getFlit)
			, .EN_recv_ports_51_putNonFullVCs(1'b1)
			, .recv_ports_51_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_51_getRecvPortID(recv_ports_info_51_getRecvPortID)
			

			, .send_ports_52_putFlit_flit_in(send_ports_52_putFlit_flit_in)
			, .EN_send_ports_52_putFlit(EN_send_ports_52_putFlit)
			, .EN_send_ports_52_getNonFullVCs(1'b1)
			, .send_ports_52_getNonFullVCs(send_ports_52_getNonFullVCs)
			, .recv_ports_52_getFlit(recv_ports_52_getFlit)
			, .EN_recv_ports_52_getFlit(EN_recv_ports_52_getFlit)
			, .EN_recv_ports_52_putNonFullVCs(1'b1)
			, .recv_ports_52_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_52_getRecvPortID(recv_ports_info_52_getRecvPortID)
			

			, .send_ports_53_putFlit_flit_in(send_ports_53_putFlit_flit_in)
			, .EN_send_ports_53_putFlit(EN_send_ports_53_putFlit)
			, .EN_send_ports_53_getNonFullVCs(1'b1)
			, .send_ports_53_getNonFullVCs(send_ports_53_getNonFullVCs)
			, .recv_ports_53_getFlit(recv_ports_53_getFlit)
			, .EN_recv_ports_53_getFlit(EN_recv_ports_53_getFlit)
			, .EN_recv_ports_53_putNonFullVCs(1'b1)
			, .recv_ports_53_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_53_getRecvPortID(recv_ports_info_53_getRecvPortID)
			

			, .send_ports_54_putFlit_flit_in(send_ports_54_putFlit_flit_in)
			, .EN_send_ports_54_putFlit(EN_send_ports_54_putFlit)
			, .EN_send_ports_54_getNonFullVCs(1'b1)
			, .send_ports_54_getNonFullVCs(send_ports_54_getNonFullVCs)
			, .recv_ports_54_getFlit(recv_ports_54_getFlit)
			, .EN_recv_ports_54_getFlit(EN_recv_ports_54_getFlit)
			, .EN_recv_ports_54_putNonFullVCs(1'b1)
			, .recv_ports_54_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_54_getRecvPortID(recv_ports_info_54_getRecvPortID)
			

			, .send_ports_55_putFlit_flit_in(send_ports_55_putFlit_flit_in)
			, .EN_send_ports_55_putFlit(EN_send_ports_55_putFlit)
			, .EN_send_ports_55_getNonFullVCs(1'b1)
			, .send_ports_55_getNonFullVCs(send_ports_55_getNonFullVCs)
			, .recv_ports_55_getFlit(recv_ports_55_getFlit)
			, .EN_recv_ports_55_getFlit(EN_recv_ports_55_getFlit)
			, .EN_recv_ports_55_putNonFullVCs(1'b1)
			, .recv_ports_55_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_55_getRecvPortID(recv_ports_info_55_getRecvPortID)
			

			, .send_ports_56_putFlit_flit_in(send_ports_56_putFlit_flit_in)
			, .EN_send_ports_56_putFlit(EN_send_ports_56_putFlit)
			, .EN_send_ports_56_getNonFullVCs(1'b1)
			, .send_ports_56_getNonFullVCs(send_ports_56_getNonFullVCs)
			, .recv_ports_56_getFlit(recv_ports_56_getFlit)
			, .EN_recv_ports_56_getFlit(EN_recv_ports_56_getFlit)
			, .EN_recv_ports_56_putNonFullVCs(1'b1)
			, .recv_ports_56_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_56_getRecvPortID(recv_ports_info_56_getRecvPortID)
			

			, .send_ports_57_putFlit_flit_in(send_ports_57_putFlit_flit_in)
			, .EN_send_ports_57_putFlit(EN_send_ports_57_putFlit)
			, .EN_send_ports_57_getNonFullVCs(1'b1)
			, .send_ports_57_getNonFullVCs(send_ports_57_getNonFullVCs)
			, .recv_ports_57_getFlit(recv_ports_57_getFlit)
			, .EN_recv_ports_57_getFlit(EN_recv_ports_57_getFlit)
			, .EN_recv_ports_57_putNonFullVCs(1'b1)
			, .recv_ports_57_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_57_getRecvPortID(recv_ports_info_57_getRecvPortID)
			

			, .send_ports_58_putFlit_flit_in(send_ports_58_putFlit_flit_in)
			, .EN_send_ports_58_putFlit(EN_send_ports_58_putFlit)
			, .EN_send_ports_58_getNonFullVCs(1'b1)
			, .send_ports_58_getNonFullVCs(send_ports_58_getNonFullVCs)
			, .recv_ports_58_getFlit(recv_ports_58_getFlit)
			, .EN_recv_ports_58_getFlit(EN_recv_ports_58_getFlit)
			, .EN_recv_ports_58_putNonFullVCs(1'b1)
			, .recv_ports_58_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_58_getRecvPortID(recv_ports_info_58_getRecvPortID)
			

			, .send_ports_59_putFlit_flit_in(send_ports_59_putFlit_flit_in)
			, .EN_send_ports_59_putFlit(EN_send_ports_59_putFlit)
			, .EN_send_ports_59_getNonFullVCs(1'b1)
			, .send_ports_59_getNonFullVCs(send_ports_59_getNonFullVCs)
			, .recv_ports_59_getFlit(recv_ports_59_getFlit)
			, .EN_recv_ports_59_getFlit(EN_recv_ports_59_getFlit)
			, .EN_recv_ports_59_putNonFullVCs(1'b1)
			, .recv_ports_59_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_59_getRecvPortID(recv_ports_info_59_getRecvPortID)
			

			, .send_ports_60_putFlit_flit_in(send_ports_60_putFlit_flit_in)
			, .EN_send_ports_60_putFlit(EN_send_ports_60_putFlit)
			, .EN_send_ports_60_getNonFullVCs(1'b1)
			, .send_ports_60_getNonFullVCs(send_ports_60_getNonFullVCs)
			, .recv_ports_60_getFlit(recv_ports_60_getFlit)
			, .EN_recv_ports_60_getFlit(EN_recv_ports_60_getFlit)
			, .EN_recv_ports_60_putNonFullVCs(1'b1)
			, .recv_ports_60_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_60_getRecvPortID(recv_ports_info_60_getRecvPortID)
			

			, .send_ports_61_putFlit_flit_in(send_ports_61_putFlit_flit_in)
			, .EN_send_ports_61_putFlit(EN_send_ports_61_putFlit)
			, .EN_send_ports_61_getNonFullVCs(1'b1)
			, .send_ports_61_getNonFullVCs(send_ports_61_getNonFullVCs)
			, .recv_ports_61_getFlit(recv_ports_61_getFlit)
			, .EN_recv_ports_61_getFlit(EN_recv_ports_61_getFlit)
			, .EN_recv_ports_61_putNonFullVCs(1'b1)
			, .recv_ports_61_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_61_getRecvPortID(recv_ports_info_61_getRecvPortID)
			

			, .send_ports_62_putFlit_flit_in(send_ports_62_putFlit_flit_in)
			, .EN_send_ports_62_putFlit(EN_send_ports_62_putFlit)
			, .EN_send_ports_62_getNonFullVCs(1'b1)
			, .send_ports_62_getNonFullVCs(send_ports_62_getNonFullVCs)
			, .recv_ports_62_getFlit(recv_ports_62_getFlit)
			, .EN_recv_ports_62_getFlit(EN_recv_ports_62_getFlit)
			, .EN_recv_ports_62_putNonFullVCs(1'b1)
			, .recv_ports_62_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_62_getRecvPortID(recv_ports_info_62_getRecvPortID)
			

			, .send_ports_63_putFlit_flit_in(send_ports_63_putFlit_flit_in)
			, .EN_send_ports_63_putFlit(EN_send_ports_63_putFlit)
			, .EN_send_ports_63_getNonFullVCs(1'b1)
			, .send_ports_63_getNonFullVCs(send_ports_63_getNonFullVCs)
			, .recv_ports_63_getFlit(recv_ports_63_getFlit)
			, .EN_recv_ports_63_getFlit(EN_recv_ports_63_getFlit)
			, .EN_recv_ports_63_putNonFullVCs(1'b1)
			, .recv_ports_63_putNonFullVCs_nonFullVCs('b1)
			, .recv_ports_info_63_getRecvPortID(recv_ports_info_63_getRecvPortID)
			

	);


	multNode node_0 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_0_getRecvPortID),
				.getVertex(getVertex_0),
				.flit_in(recv_ports_0_getFlit),
				.rcvReady(EN_recv_ports_0_getFlit),
				.canSend(send_ports_0_getNonFullVCs[0]),
				.flit_out(send_ports_0_putFlit_flit_in),
				.putFlit(EN_send_ports_0_putFlit),
				.LUT_address(LUT_address_0),
				.LUT_output_data(LUT_output_data_0),
				.vertex(vertex_0),
				.done(done)
		);

 
	multNode node_1 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_1_getRecvPortID),
				.getVertex(getVertex_1),
				.flit_in(recv_ports_1_getFlit),
				.rcvReady(EN_recv_ports_1_getFlit),
				.canSend(send_ports_1_getNonFullVCs[0]),
				.flit_out(send_ports_1_putFlit_flit_in),
				.putFlit(EN_send_ports_1_putFlit),
				.LUT_address(LUT_address_1),
				.LUT_output_data(LUT_output_data_1),
				.vertex(vertex_1)
		);

 
	multNode node_2 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_2_getRecvPortID),
				.getVertex(getVertex_2),
				.flit_in(recv_ports_2_getFlit),
				.rcvReady(EN_recv_ports_2_getFlit),
				.canSend(send_ports_2_getNonFullVCs[0]),
				.flit_out(send_ports_2_putFlit_flit_in),
				.putFlit(EN_send_ports_2_putFlit),
				.LUT_address(LUT_address_2),
				.LUT_output_data(LUT_output_data_2),
				.vertex(vertex_2)
		);

 
	multNode node_3 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_3_getRecvPortID),
				.getVertex(getVertex_3),
				.flit_in(recv_ports_3_getFlit),
				.rcvReady(EN_recv_ports_3_getFlit),
				.canSend(send_ports_3_getNonFullVCs[0]),
				.flit_out(send_ports_3_putFlit_flit_in),
				.putFlit(EN_send_ports_3_putFlit),
				.LUT_address(LUT_address_3),
				.LUT_output_data(LUT_output_data_3),
				.vertex(vertex_3)
		);

 
	multNode node_4 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_4_getRecvPortID),
				.getVertex(getVertex_4),
				.flit_in(recv_ports_4_getFlit),
				.rcvReady(EN_recv_ports_4_getFlit),
				.canSend(send_ports_4_getNonFullVCs[0]),
				.flit_out(send_ports_4_putFlit_flit_in),
				.putFlit(EN_send_ports_4_putFlit),
				.LUT_address(LUT_address_4),
				.LUT_output_data(LUT_output_data_4),
				.vertex(vertex_4)
		);

 
	multNode node_5 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_5_getRecvPortID),
				.getVertex(getVertex_5),
				.flit_in(recv_ports_5_getFlit),
				.rcvReady(EN_recv_ports_5_getFlit),
				.canSend(send_ports_5_getNonFullVCs[0]),
				.flit_out(send_ports_5_putFlit_flit_in),
				.putFlit(EN_send_ports_5_putFlit),
				.LUT_address(LUT_address_5),
				.LUT_output_data(LUT_output_data_5),
				.vertex(vertex_5)
		);

 
	multNode node_6 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_6_getRecvPortID),
				.getVertex(getVertex_6),
				.flit_in(recv_ports_6_getFlit),
				.rcvReady(EN_recv_ports_6_getFlit),
				.canSend(send_ports_6_getNonFullVCs[0]),
				.flit_out(send_ports_6_putFlit_flit_in),
				.putFlit(EN_send_ports_6_putFlit),
				.LUT_address(LUT_address_6),
				.LUT_output_data(LUT_output_data_6),
				.vertex(vertex_6)
		);

 
	multNode node_7 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_7_getRecvPortID),
				.getVertex(getVertex_7),
				.flit_in(recv_ports_7_getFlit),
				.rcvReady(EN_recv_ports_7_getFlit),
				.canSend(send_ports_7_getNonFullVCs[0]),
				.flit_out(send_ports_7_putFlit_flit_in),
				.putFlit(EN_send_ports_7_putFlit),
				.LUT_address(LUT_address_7),
				.LUT_output_data(LUT_output_data_7),
				.vertex(vertex_7)
		);

 
	multNode node_8 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_8_getRecvPortID),
				.getVertex(getVertex_8),
				.flit_in(recv_ports_8_getFlit),
				.rcvReady(EN_recv_ports_8_getFlit),
				.canSend(send_ports_8_getNonFullVCs[0]),
				.flit_out(send_ports_8_putFlit_flit_in),
				.putFlit(EN_send_ports_8_putFlit),
				.LUT_address(LUT_address_8),
				.LUT_output_data(LUT_output_data_8),
				.vertex(vertex_8)
		);

 
	multNode node_9 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_9_getRecvPortID),
				.getVertex(getVertex_9),
				.flit_in(recv_ports_9_getFlit),
				.rcvReady(EN_recv_ports_9_getFlit),
				.canSend(send_ports_9_getNonFullVCs[0]),
				.flit_out(send_ports_9_putFlit_flit_in),
				.putFlit(EN_send_ports_9_putFlit),
				.LUT_address(LUT_address_9),
				.LUT_output_data(LUT_output_data_9),
				.vertex(vertex_9)
		);

 
	multNode node_10 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_10_getRecvPortID),
				.getVertex(getVertex_10),
				.flit_in(recv_ports_10_getFlit),
				.rcvReady(EN_recv_ports_10_getFlit),
				.canSend(send_ports_10_getNonFullVCs[0]),
				.flit_out(send_ports_10_putFlit_flit_in),
				.putFlit(EN_send_ports_10_putFlit),
				.LUT_address(LUT_address_10),
				.LUT_output_data(LUT_output_data_10),
				.vertex(vertex_10)
		);

 
	multNode node_11 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_11_getRecvPortID),
				.getVertex(getVertex_11),
				.flit_in(recv_ports_11_getFlit),
				.rcvReady(EN_recv_ports_11_getFlit),
				.canSend(send_ports_11_getNonFullVCs[0]),
				.flit_out(send_ports_11_putFlit_flit_in),
				.putFlit(EN_send_ports_11_putFlit),
				.LUT_address(LUT_address_11),
				.LUT_output_data(LUT_output_data_11),
				.vertex(vertex_11)
		);

 
	multNode node_12 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_12_getRecvPortID),
				.getVertex(getVertex_12),
				.flit_in(recv_ports_12_getFlit),
				.rcvReady(EN_recv_ports_12_getFlit),
				.canSend(send_ports_12_getNonFullVCs[0]),
				.flit_out(send_ports_12_putFlit_flit_in),
				.putFlit(EN_send_ports_12_putFlit),
				.LUT_address(LUT_address_12),
				.LUT_output_data(LUT_output_data_12),
				.vertex(vertex_12)
		);

 
	multNode node_13 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_13_getRecvPortID),
				.getVertex(getVertex_13),
				.flit_in(recv_ports_13_getFlit),
				.rcvReady(EN_recv_ports_13_getFlit),
				.canSend(send_ports_13_getNonFullVCs[0]),
				.flit_out(send_ports_13_putFlit_flit_in),
				.putFlit(EN_send_ports_13_putFlit),
				.LUT_address(LUT_address_13),
				.LUT_output_data(LUT_output_data_13),
				.vertex(vertex_13)
		);

 
	multNode node_14 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_14_getRecvPortID),
				.getVertex(getVertex_14),
				.flit_in(recv_ports_14_getFlit),
				.rcvReady(EN_recv_ports_14_getFlit),
				.canSend(send_ports_14_getNonFullVCs[0]),
				.flit_out(send_ports_14_putFlit_flit_in),
				.putFlit(EN_send_ports_14_putFlit),
				.LUT_address(LUT_address_14),
				.LUT_output_data(LUT_output_data_14),
				.vertex(vertex_14)
		);

 
	multNode node_15 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_15_getRecvPortID),
				.getVertex(getVertex_15),
				.flit_in(recv_ports_15_getFlit),
				.rcvReady(EN_recv_ports_15_getFlit),
				.canSend(send_ports_15_getNonFullVCs[0]),
				.flit_out(send_ports_15_putFlit_flit_in),
				.putFlit(EN_send_ports_15_putFlit),
				.LUT_address(LUT_address_15),
				.LUT_output_data(LUT_output_data_15),
				.vertex(vertex_15)
		);

 
	multNode node_16 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_16_getRecvPortID),
				.getVertex(getVertex_16),
				.flit_in(recv_ports_16_getFlit),
				.rcvReady(EN_recv_ports_16_getFlit),
				.canSend(send_ports_16_getNonFullVCs[0]),
				.flit_out(send_ports_16_putFlit_flit_in),
				.putFlit(EN_send_ports_16_putFlit),
				.LUT_address(LUT_address_16),
				.LUT_output_data(LUT_output_data_16),
				.vertex(vertex_16)
		);

 
	multNode node_17 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_17_getRecvPortID),
				.getVertex(getVertex_17),
				.flit_in(recv_ports_17_getFlit),
				.rcvReady(EN_recv_ports_17_getFlit),
				.canSend(send_ports_17_getNonFullVCs[0]),
				.flit_out(send_ports_17_putFlit_flit_in),
				.putFlit(EN_send_ports_17_putFlit),
				.LUT_address(LUT_address_17),
				.LUT_output_data(LUT_output_data_17),
				.vertex(vertex_17)
		);

 
	multNode node_18 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_18_getRecvPortID),
				.getVertex(getVertex_18),
				.flit_in(recv_ports_18_getFlit),
				.rcvReady(EN_recv_ports_18_getFlit),
				.canSend(send_ports_18_getNonFullVCs[0]),
				.flit_out(send_ports_18_putFlit_flit_in),
				.putFlit(EN_send_ports_18_putFlit),
				.LUT_address(LUT_address_18),
				.LUT_output_data(LUT_output_data_18),
				.vertex(vertex_18)
		);

 
	multNode node_19 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_19_getRecvPortID),
				.getVertex(getVertex_19),
				.flit_in(recv_ports_19_getFlit),
				.rcvReady(EN_recv_ports_19_getFlit),
				.canSend(send_ports_19_getNonFullVCs[0]),
				.flit_out(send_ports_19_putFlit_flit_in),
				.putFlit(EN_send_ports_19_putFlit),
				.LUT_address(LUT_address_19),
				.LUT_output_data(LUT_output_data_19),
				.vertex(vertex_19)
		);

 
	multNode node_20 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_20_getRecvPortID),
				.getVertex(getVertex_20),
				.flit_in(recv_ports_20_getFlit),
				.rcvReady(EN_recv_ports_20_getFlit),
				.canSend(send_ports_20_getNonFullVCs[0]),
				.flit_out(send_ports_20_putFlit_flit_in),
				.putFlit(EN_send_ports_20_putFlit),
				.LUT_address(LUT_address_20),
				.LUT_output_data(LUT_output_data_20),
				.vertex(vertex_20)
		);

 
	multNode node_21 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_21_getRecvPortID),
				.getVertex(getVertex_21),
				.flit_in(recv_ports_21_getFlit),
				.rcvReady(EN_recv_ports_21_getFlit),
				.canSend(send_ports_21_getNonFullVCs[0]),
				.flit_out(send_ports_21_putFlit_flit_in),
				.putFlit(EN_send_ports_21_putFlit),
				.LUT_address(LUT_address_21),
				.LUT_output_data(LUT_output_data_21),
				.vertex(vertex_21)
		);

 
	multNode node_22 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_22_getRecvPortID),
				.getVertex(getVertex_22),
				.flit_in(recv_ports_22_getFlit),
				.rcvReady(EN_recv_ports_22_getFlit),
				.canSend(send_ports_22_getNonFullVCs[0]),
				.flit_out(send_ports_22_putFlit_flit_in),
				.putFlit(EN_send_ports_22_putFlit),
				.LUT_address(LUT_address_22),
				.LUT_output_data(LUT_output_data_22),
				.vertex(vertex_22)
		);

 
	multNode node_23 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_23_getRecvPortID),
				.getVertex(getVertex_23),
				.flit_in(recv_ports_23_getFlit),
				.rcvReady(EN_recv_ports_23_getFlit),
				.canSend(send_ports_23_getNonFullVCs[0]),
				.flit_out(send_ports_23_putFlit_flit_in),
				.putFlit(EN_send_ports_23_putFlit),
				.LUT_address(LUT_address_23),
				.LUT_output_data(LUT_output_data_23),
				.vertex(vertex_23)
		);

 
	multNode node_24 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_24_getRecvPortID),
				.getVertex(getVertex_24),
				.flit_in(recv_ports_24_getFlit),
				.rcvReady(EN_recv_ports_24_getFlit),
				.canSend(send_ports_24_getNonFullVCs[0]),
				.flit_out(send_ports_24_putFlit_flit_in),
				.putFlit(EN_send_ports_24_putFlit),
				.LUT_address(LUT_address_24),
				.LUT_output_data(LUT_output_data_24),
				.vertex(vertex_24)
		);

 
	multNode node_25 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_25_getRecvPortID),
				.getVertex(getVertex_25),
				.flit_in(recv_ports_25_getFlit),
				.rcvReady(EN_recv_ports_25_getFlit),
				.canSend(send_ports_25_getNonFullVCs[0]),
				.flit_out(send_ports_25_putFlit_flit_in),
				.putFlit(EN_send_ports_25_putFlit),
				.LUT_address(LUT_address_25),
				.LUT_output_data(LUT_output_data_25),
				.vertex(vertex_25)
		);

 
	multNode node_26 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_26_getRecvPortID),
				.getVertex(getVertex_26),
				.flit_in(recv_ports_26_getFlit),
				.rcvReady(EN_recv_ports_26_getFlit),
				.canSend(send_ports_26_getNonFullVCs[0]),
				.flit_out(send_ports_26_putFlit_flit_in),
				.putFlit(EN_send_ports_26_putFlit),
				.LUT_address(LUT_address_26),
				.LUT_output_data(LUT_output_data_26),
				.vertex(vertex_26)
		);

 
	multNode node_27 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_27_getRecvPortID),
				.getVertex(getVertex_27),
				.flit_in(recv_ports_27_getFlit),
				.rcvReady(EN_recv_ports_27_getFlit),
				.canSend(send_ports_27_getNonFullVCs[0]),
				.flit_out(send_ports_27_putFlit_flit_in),
				.putFlit(EN_send_ports_27_putFlit),
				.LUT_address(LUT_address_27),
				.LUT_output_data(LUT_output_data_27),
				.vertex(vertex_27)
		);

 
	multNode node_28 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_28_getRecvPortID),
				.getVertex(getVertex_28),
				.flit_in(recv_ports_28_getFlit),
				.rcvReady(EN_recv_ports_28_getFlit),
				.canSend(send_ports_28_getNonFullVCs[0]),
				.flit_out(send_ports_28_putFlit_flit_in),
				.putFlit(EN_send_ports_28_putFlit),
				.LUT_address(LUT_address_28),
				.LUT_output_data(LUT_output_data_28),
				.vertex(vertex_28)
		);

 
	multNode node_29 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_29_getRecvPortID),
				.getVertex(getVertex_29),
				.flit_in(recv_ports_29_getFlit),
				.rcvReady(EN_recv_ports_29_getFlit),
				.canSend(send_ports_29_getNonFullVCs[0]),
				.flit_out(send_ports_29_putFlit_flit_in),
				.putFlit(EN_send_ports_29_putFlit),
				.LUT_address(LUT_address_29),
				.LUT_output_data(LUT_output_data_29),
				.vertex(vertex_29)
		);

 
	multNode node_30 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_30_getRecvPortID),
				.getVertex(getVertex_30),
				.flit_in(recv_ports_30_getFlit),
				.rcvReady(EN_recv_ports_30_getFlit),
				.canSend(send_ports_30_getNonFullVCs[0]),
				.flit_out(send_ports_30_putFlit_flit_in),
				.putFlit(EN_send_ports_30_putFlit),
				.LUT_address(LUT_address_30),
				.LUT_output_data(LUT_output_data_30),
				.vertex(vertex_30)
		);

 
	multNode node_31 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_31_getRecvPortID),
				.getVertex(getVertex_31),
				.flit_in(recv_ports_31_getFlit),
				.rcvReady(EN_recv_ports_31_getFlit),
				.canSend(send_ports_31_getNonFullVCs[0]),
				.flit_out(send_ports_31_putFlit_flit_in),
				.putFlit(EN_send_ports_31_putFlit),
				.LUT_address(LUT_address_31),
				.LUT_output_data(LUT_output_data_31),
				.vertex(vertex_31)
		);

 
	multNode node_32 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_32_getRecvPortID),
				.getVertex(getVertex_32),
				.flit_in(recv_ports_32_getFlit),
				.rcvReady(EN_recv_ports_32_getFlit),
				.canSend(send_ports_32_getNonFullVCs[0]),
				.flit_out(send_ports_32_putFlit_flit_in),
				.putFlit(EN_send_ports_32_putFlit),
				.LUT_address(LUT_address_32),
				.LUT_output_data(LUT_output_data_32),
				.vertex(vertex_32)
		);

 
	multNode node_33 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_33_getRecvPortID),
				.getVertex(getVertex_33),
				.flit_in(recv_ports_33_getFlit),
				.rcvReady(EN_recv_ports_33_getFlit),
				.canSend(send_ports_33_getNonFullVCs[0]),
				.flit_out(send_ports_33_putFlit_flit_in),
				.putFlit(EN_send_ports_33_putFlit),
				.LUT_address(LUT_address_33),
				.LUT_output_data(LUT_output_data_33),
				.vertex(vertex_33)
		);

 
	multNode node_34 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_34_getRecvPortID),
				.getVertex(getVertex_34),
				.flit_in(recv_ports_34_getFlit),
				.rcvReady(EN_recv_ports_34_getFlit),
				.canSend(send_ports_34_getNonFullVCs[0]),
				.flit_out(send_ports_34_putFlit_flit_in),
				.putFlit(EN_send_ports_34_putFlit),
				.LUT_address(LUT_address_34),
				.LUT_output_data(LUT_output_data_34),
				.vertex(vertex_34)
		);

 
	multNode node_35 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_35_getRecvPortID),
				.getVertex(getVertex_35),
				.flit_in(recv_ports_35_getFlit),
				.rcvReady(EN_recv_ports_35_getFlit),
				.canSend(send_ports_35_getNonFullVCs[0]),
				.flit_out(send_ports_35_putFlit_flit_in),
				.putFlit(EN_send_ports_35_putFlit),
				.LUT_address(LUT_address_35),
				.LUT_output_data(LUT_output_data_35),
				.vertex(vertex_35)
		);

 
	multNode node_36 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_36_getRecvPortID),
				.getVertex(getVertex_36),
				.flit_in(recv_ports_36_getFlit),
				.rcvReady(EN_recv_ports_36_getFlit),
				.canSend(send_ports_36_getNonFullVCs[0]),
				.flit_out(send_ports_36_putFlit_flit_in),
				.putFlit(EN_send_ports_36_putFlit),
				.LUT_address(LUT_address_36),
				.LUT_output_data(LUT_output_data_36),
				.vertex(vertex_36)
		);

 
	multNode node_37 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_37_getRecvPortID),
				.getVertex(getVertex_37),
				.flit_in(recv_ports_37_getFlit),
				.rcvReady(EN_recv_ports_37_getFlit),
				.canSend(send_ports_37_getNonFullVCs[0]),
				.flit_out(send_ports_37_putFlit_flit_in),
				.putFlit(EN_send_ports_37_putFlit),
				.LUT_address(LUT_address_37),
				.LUT_output_data(LUT_output_data_37),
				.vertex(vertex_37)
		);

 
	multNode node_38 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_38_getRecvPortID),
				.getVertex(getVertex_38),
				.flit_in(recv_ports_38_getFlit),
				.rcvReady(EN_recv_ports_38_getFlit),
				.canSend(send_ports_38_getNonFullVCs[0]),
				.flit_out(send_ports_38_putFlit_flit_in),
				.putFlit(EN_send_ports_38_putFlit),
				.LUT_address(LUT_address_38),
				.LUT_output_data(LUT_output_data_38),
				.vertex(vertex_38)
		);

 
	multNode node_39 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_39_getRecvPortID),
				.getVertex(getVertex_39),
				.flit_in(recv_ports_39_getFlit),
				.rcvReady(EN_recv_ports_39_getFlit),
				.canSend(send_ports_39_getNonFullVCs[0]),
				.flit_out(send_ports_39_putFlit_flit_in),
				.putFlit(EN_send_ports_39_putFlit),
				.LUT_address(LUT_address_39),
				.LUT_output_data(LUT_output_data_39),
				.vertex(vertex_39)
		);

 
	multNode node_40 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_40_getRecvPortID),
				.getVertex(getVertex_40),
				.flit_in(recv_ports_40_getFlit),
				.rcvReady(EN_recv_ports_40_getFlit),
				.canSend(send_ports_40_getNonFullVCs[0]),
				.flit_out(send_ports_40_putFlit_flit_in),
				.putFlit(EN_send_ports_40_putFlit),
				.LUT_address(LUT_address_40),
				.LUT_output_data(LUT_output_data_40),
				.vertex(vertex_40)
		);

 
	multNode node_41 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_41_getRecvPortID),
				.getVertex(getVertex_41),
				.flit_in(recv_ports_41_getFlit),
				.rcvReady(EN_recv_ports_41_getFlit),
				.canSend(send_ports_41_getNonFullVCs[0]),
				.flit_out(send_ports_41_putFlit_flit_in),
				.putFlit(EN_send_ports_41_putFlit),
				.LUT_address(LUT_address_41),
				.LUT_output_data(LUT_output_data_41),
				.vertex(vertex_41)
		);

 
	multNode node_42 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_42_getRecvPortID),
				.getVertex(getVertex_42),
				.flit_in(recv_ports_42_getFlit),
				.rcvReady(EN_recv_ports_42_getFlit),
				.canSend(send_ports_42_getNonFullVCs[0]),
				.flit_out(send_ports_42_putFlit_flit_in),
				.putFlit(EN_send_ports_42_putFlit),
				.LUT_address(LUT_address_42),
				.LUT_output_data(LUT_output_data_42),
				.vertex(vertex_42)
		);

 
	multNode node_43 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_43_getRecvPortID),
				.getVertex(getVertex_43),
				.flit_in(recv_ports_43_getFlit),
				.rcvReady(EN_recv_ports_43_getFlit),
				.canSend(send_ports_43_getNonFullVCs[0]),
				.flit_out(send_ports_43_putFlit_flit_in),
				.putFlit(EN_send_ports_43_putFlit),
				.LUT_address(LUT_address_43),
				.LUT_output_data(LUT_output_data_43),
				.vertex(vertex_43)
		);

 
	multNode node_44 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_44_getRecvPortID),
				.getVertex(getVertex_44),
				.flit_in(recv_ports_44_getFlit),
				.rcvReady(EN_recv_ports_44_getFlit),
				.canSend(send_ports_44_getNonFullVCs[0]),
				.flit_out(send_ports_44_putFlit_flit_in),
				.putFlit(EN_send_ports_44_putFlit),
				.LUT_address(LUT_address_44),
				.LUT_output_data(LUT_output_data_44),
				.vertex(vertex_44)
		);

 
	multNode node_45 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_45_getRecvPortID),
				.getVertex(getVertex_45),
				.flit_in(recv_ports_45_getFlit),
				.rcvReady(EN_recv_ports_45_getFlit),
				.canSend(send_ports_45_getNonFullVCs[0]),
				.flit_out(send_ports_45_putFlit_flit_in),
				.putFlit(EN_send_ports_45_putFlit),
				.LUT_address(LUT_address_45),
				.LUT_output_data(LUT_output_data_45),
				.vertex(vertex_45)
		);

 
	multNode node_46 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_46_getRecvPortID),
				.getVertex(getVertex_46),
				.flit_in(recv_ports_46_getFlit),
				.rcvReady(EN_recv_ports_46_getFlit),
				.canSend(send_ports_46_getNonFullVCs[0]),
				.flit_out(send_ports_46_putFlit_flit_in),
				.putFlit(EN_send_ports_46_putFlit),
				.LUT_address(LUT_address_46),
				.LUT_output_data(LUT_output_data_46),
				.vertex(vertex_46)
		);

 
	multNode node_47 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_47_getRecvPortID),
				.getVertex(getVertex_47),
				.flit_in(recv_ports_47_getFlit),
				.rcvReady(EN_recv_ports_47_getFlit),
				.canSend(send_ports_47_getNonFullVCs[0]),
				.flit_out(send_ports_47_putFlit_flit_in),
				.putFlit(EN_send_ports_47_putFlit),
				.LUT_address(LUT_address_47),
				.LUT_output_data(LUT_output_data_47),
				.vertex(vertex_47)
		);

 
	multNode node_48 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_48_getRecvPortID),
				.getVertex(getVertex_48),
				.flit_in(recv_ports_48_getFlit),
				.rcvReady(EN_recv_ports_48_getFlit),
				.canSend(send_ports_48_getNonFullVCs[0]),
				.flit_out(send_ports_48_putFlit_flit_in),
				.putFlit(EN_send_ports_48_putFlit),
				.LUT_address(LUT_address_48),
				.LUT_output_data(LUT_output_data_48),
				.vertex(vertex_48)
		);

 
	multNode node_49 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_49_getRecvPortID),
				.getVertex(getVertex_49),
				.flit_in(recv_ports_49_getFlit),
				.rcvReady(EN_recv_ports_49_getFlit),
				.canSend(send_ports_49_getNonFullVCs[0]),
				.flit_out(send_ports_49_putFlit_flit_in),
				.putFlit(EN_send_ports_49_putFlit),
				.LUT_address(LUT_address_49),
				.LUT_output_data(LUT_output_data_49),
				.vertex(vertex_49)
		);

 
	multNode node_50 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_50_getRecvPortID),
				.getVertex(getVertex_50),
				.flit_in(recv_ports_50_getFlit),
				.rcvReady(EN_recv_ports_50_getFlit),
				.canSend(send_ports_50_getNonFullVCs[0]),
				.flit_out(send_ports_50_putFlit_flit_in),
				.putFlit(EN_send_ports_50_putFlit),
				.LUT_address(LUT_address_50),
				.LUT_output_data(LUT_output_data_50),
				.vertex(vertex_50)
		);

 
	multNode node_51 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_51_getRecvPortID),
				.getVertex(getVertex_51),
				.flit_in(recv_ports_51_getFlit),
				.rcvReady(EN_recv_ports_51_getFlit),
				.canSend(send_ports_51_getNonFullVCs[0]),
				.flit_out(send_ports_51_putFlit_flit_in),
				.putFlit(EN_send_ports_51_putFlit),
				.LUT_address(LUT_address_51),
				.LUT_output_data(LUT_output_data_51),
				.vertex(vertex_51)
		);

 
	multNode node_52 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_52_getRecvPortID),
				.getVertex(getVertex_52),
				.flit_in(recv_ports_52_getFlit),
				.rcvReady(EN_recv_ports_52_getFlit),
				.canSend(send_ports_52_getNonFullVCs[0]),
				.flit_out(send_ports_52_putFlit_flit_in),
				.putFlit(EN_send_ports_52_putFlit),
				.LUT_address(LUT_address_52),
				.LUT_output_data(LUT_output_data_52),
				.vertex(vertex_52)
		);

 
	multNode node_53 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_53_getRecvPortID),
				.getVertex(getVertex_53),
				.flit_in(recv_ports_53_getFlit),
				.rcvReady(EN_recv_ports_53_getFlit),
				.canSend(send_ports_53_getNonFullVCs[0]),
				.flit_out(send_ports_53_putFlit_flit_in),
				.putFlit(EN_send_ports_53_putFlit),
				.LUT_address(LUT_address_53),
				.LUT_output_data(LUT_output_data_53),
				.vertex(vertex_53)
		);

 
	multNode node_54 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_54_getRecvPortID),
				.getVertex(getVertex_54),
				.flit_in(recv_ports_54_getFlit),
				.rcvReady(EN_recv_ports_54_getFlit),
				.canSend(send_ports_54_getNonFullVCs[0]),
				.flit_out(send_ports_54_putFlit_flit_in),
				.putFlit(EN_send_ports_54_putFlit),
				.LUT_address(LUT_address_54),
				.LUT_output_data(LUT_output_data_54),
				.vertex(vertex_54)
		);

 
	multNode node_55 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_55_getRecvPortID),
				.getVertex(getVertex_55),
				.flit_in(recv_ports_55_getFlit),
				.rcvReady(EN_recv_ports_55_getFlit),
				.canSend(send_ports_55_getNonFullVCs[0]),
				.flit_out(send_ports_55_putFlit_flit_in),
				.putFlit(EN_send_ports_55_putFlit),
				.LUT_address(LUT_address_55),
				.LUT_output_data(LUT_output_data_55),
				.vertex(vertex_55)
		);

 
	multNode node_56 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_56_getRecvPortID),
				.getVertex(getVertex_56),
				.flit_in(recv_ports_56_getFlit),
				.rcvReady(EN_recv_ports_56_getFlit),
				.canSend(send_ports_56_getNonFullVCs[0]),
				.flit_out(send_ports_56_putFlit_flit_in),
				.putFlit(EN_send_ports_56_putFlit),
				.LUT_address(LUT_address_56),
				.LUT_output_data(LUT_output_data_56),
				.vertex(vertex_56)
		);

 
	multNode node_57 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_57_getRecvPortID),
				.getVertex(getVertex_57),
				.flit_in(recv_ports_57_getFlit),
				.rcvReady(EN_recv_ports_57_getFlit),
				.canSend(send_ports_57_getNonFullVCs[0]),
				.flit_out(send_ports_57_putFlit_flit_in),
				.putFlit(EN_send_ports_57_putFlit),
				.LUT_address(LUT_address_57),
				.LUT_output_data(LUT_output_data_57),
				.vertex(vertex_57)
		);

 
	multNode node_58 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_58_getRecvPortID),
				.getVertex(getVertex_58),
				.flit_in(recv_ports_58_getFlit),
				.rcvReady(EN_recv_ports_58_getFlit),
				.canSend(send_ports_58_getNonFullVCs[0]),
				.flit_out(send_ports_58_putFlit_flit_in),
				.putFlit(EN_send_ports_58_putFlit),
				.LUT_address(LUT_address_58),
				.LUT_output_data(LUT_output_data_58),
				.vertex(vertex_58)
		);

 
	multNode node_59 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_59_getRecvPortID),
				.getVertex(getVertex_59),
				.flit_in(recv_ports_59_getFlit),
				.rcvReady(EN_recv_ports_59_getFlit),
				.canSend(send_ports_59_getNonFullVCs[0]),
				.flit_out(send_ports_59_putFlit_flit_in),
				.putFlit(EN_send_ports_59_putFlit),
				.LUT_address(LUT_address_59),
				.LUT_output_data(LUT_output_data_59),
				.vertex(vertex_59)
		);

 
	multNode node_60 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_60_getRecvPortID),
				.getVertex(getVertex_60),
				.flit_in(recv_ports_60_getFlit),
				.rcvReady(EN_recv_ports_60_getFlit),
				.canSend(send_ports_60_getNonFullVCs[0]),
				.flit_out(send_ports_60_putFlit_flit_in),
				.putFlit(EN_send_ports_60_putFlit),
				.LUT_address(LUT_address_60),
				.LUT_output_data(LUT_output_data_60),
				.vertex(vertex_60)
		);

 
	multNode node_61 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_61_getRecvPortID),
				.getVertex(getVertex_61),
				.flit_in(recv_ports_61_getFlit),
				.rcvReady(EN_recv_ports_61_getFlit),
				.canSend(send_ports_61_getNonFullVCs[0]),
				.flit_out(send_ports_61_putFlit_flit_in),
				.putFlit(EN_send_ports_61_putFlit),
				.LUT_address(LUT_address_61),
				.LUT_output_data(LUT_output_data_61),
				.vertex(vertex_61)
		);

 
	multNode node_62 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_62_getRecvPortID),
				.getVertex(getVertex_62),
				.flit_in(recv_ports_62_getFlit),
				.rcvReady(EN_recv_ports_62_getFlit),
				.canSend(send_ports_62_getNonFullVCs[0]),
				.flit_out(send_ports_62_putFlit_flit_in),
				.putFlit(EN_send_ports_62_putFlit),
				.LUT_address(LUT_address_62),
				.LUT_output_data(LUT_output_data_62),
				.vertex(vertex_62)
		);

 
	multNode node_63 (
				.reset(reset),
				.clk(clk),
				.max_iteration(max_iteration),
				.getID(recv_ports_info_63_getRecvPortID),
				.getVertex(getVertex_63),
				.flit_in(recv_ports_63_getFlit),
				.rcvReady(EN_recv_ports_63_getFlit),
				.canSend(send_ports_63_getNonFullVCs[0]),
				.flit_out(send_ports_63_putFlit_flit_in),
				.putFlit(EN_send_ports_63_putFlit),
				.LUT_address(LUT_address_63),
				.LUT_output_data(LUT_output_data_63),
				.vertex(vertex_63)
		);
		
		
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_1.data") LUT_0( .clk(clk), .write_enable(1'b0), .address(LUT_address_0), .output_data(LUT_output_data_0)); 		
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_2.data") LUT_1( .clk(clk), .write_enable(1'b0), .address(LUT_address_1), .output_data(LUT_output_data_1)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_3.data") LUT_2( .clk(clk), .write_enable(1'b0), .address(LUT_address_2), .output_data(LUT_output_data_2)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_4.data") LUT_3( .clk(clk), .write_enable(1'b0), .address(LUT_address_3), .output_data(LUT_output_data_3)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_5.data") LUT_4( .clk(clk), .write_enable(1'b0), .address(LUT_address_4), .output_data(LUT_output_data_4)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_6.data") LUT_5( .clk(clk), .write_enable(1'b0), .address(LUT_address_5), .output_data(LUT_output_data_5)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_7.data") LUT_6( .clk(clk), .write_enable(1'b0), .address(LUT_address_6), .output_data(LUT_output_data_6)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_8.data") LUT_7( .clk(clk), .write_enable(1'b0), .address(LUT_address_7), .output_data(LUT_output_data_7)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_9.data") LUT_8( .clk(clk), .write_enable(1'b0), .address(LUT_address_8), .output_data(LUT_output_data_8)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_10.data") LUT_9( .clk(clk), .write_enable(1'b0), .address(LUT_address_9), .output_data(LUT_output_data_9)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_11.data") LUT_10( .clk(clk), .write_enable(1'b0), .address(LUT_address_10), .output_data(LUT_output_data_10)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_12.data") LUT_11( .clk(clk), .write_enable(1'b0), .address(LUT_address_11), .output_data(LUT_output_data_11)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_13.data") LUT_12( .clk(clk), .write_enable(1'b0), .address(LUT_address_12), .output_data(LUT_output_data_12)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_14.data") LUT_13( .clk(clk), .write_enable(1'b0), .address(LUT_address_13), .output_data(LUT_output_data_13)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_15.data") LUT_14( .clk(clk), .write_enable(1'b0), .address(LUT_address_14), .output_data(LUT_output_data_14)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_16.data") LUT_15( .clk(clk), .write_enable(1'b0), .address(LUT_address_15), .output_data(LUT_output_data_15)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_17.data") LUT_16( .clk(clk), .write_enable(1'b0), .address(LUT_address_16), .output_data(LUT_output_data_16)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_18.data") LUT_17( .clk(clk), .write_enable(1'b0), .address(LUT_address_17), .output_data(LUT_output_data_17)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_19.data") LUT_18( .clk(clk), .write_enable(1'b0), .address(LUT_address_18), .output_data(LUT_output_data_18)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_20.data") LUT_19( .clk(clk), .write_enable(1'b0), .address(LUT_address_19), .output_data(LUT_output_data_19)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_21.data") LUT_20( .clk(clk), .write_enable(1'b0), .address(LUT_address_20), .output_data(LUT_output_data_20)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_22.data") LUT_21( .clk(clk), .write_enable(1'b0), .address(LUT_address_21), .output_data(LUT_output_data_21)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_23.data") LUT_22( .clk(clk), .write_enable(1'b0), .address(LUT_address_22), .output_data(LUT_output_data_22)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_24.data") LUT_23( .clk(clk), .write_enable(1'b0), .address(LUT_address_23), .output_data(LUT_output_data_23)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_25.data") LUT_24( .clk(clk), .write_enable(1'b0), .address(LUT_address_24), .output_data(LUT_output_data_24)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_26.data") LUT_25( .clk(clk), .write_enable(1'b0), .address(LUT_address_25), .output_data(LUT_output_data_25)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_27.data") LUT_26( .clk(clk), .write_enable(1'b0), .address(LUT_address_26), .output_data(LUT_output_data_26)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_28.data") LUT_27( .clk(clk), .write_enable(1'b0), .address(LUT_address_27), .output_data(LUT_output_data_27)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_29.data") LUT_28( .clk(clk), .write_enable(1'b0), .address(LUT_address_28), .output_data(LUT_output_data_28)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_30.data") LUT_29( .clk(clk), .write_enable(1'b0), .address(LUT_address_29), .output_data(LUT_output_data_29)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_31.data") LUT_30( .clk(clk), .write_enable(1'b0), .address(LUT_address_30), .output_data(LUT_output_data_30)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_32.data") LUT_31( .clk(clk), .write_enable(1'b0), .address(LUT_address_31), .output_data(LUT_output_data_31)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_33.data") LUT_32( .clk(clk), .write_enable(1'b0), .address(LUT_address_32), .output_data(LUT_output_data_32)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_34.data") LUT_33( .clk(clk), .write_enable(1'b0), .address(LUT_address_33), .output_data(LUT_output_data_33)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_35.data") LUT_34( .clk(clk), .write_enable(1'b0), .address(LUT_address_34), .output_data(LUT_output_data_34)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_36.data") LUT_35( .clk(clk), .write_enable(1'b0), .address(LUT_address_35), .output_data(LUT_output_data_35)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_37.data") LUT_36( .clk(clk), .write_enable(1'b0), .address(LUT_address_36), .output_data(LUT_output_data_36)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_38.data") LUT_37( .clk(clk), .write_enable(1'b0), .address(LUT_address_37), .output_data(LUT_output_data_37)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_39.data") LUT_38( .clk(clk), .write_enable(1'b0), .address(LUT_address_38), .output_data(LUT_output_data_38)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_40.data") LUT_39( .clk(clk), .write_enable(1'b0), .address(LUT_address_39), .output_data(LUT_output_data_39)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_41.data") LUT_40( .clk(clk), .write_enable(1'b0), .address(LUT_address_40), .output_data(LUT_output_data_40)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_42.data") LUT_41( .clk(clk), .write_enable(1'b0), .address(LUT_address_41), .output_data(LUT_output_data_41)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_43.data") LUT_42( .clk(clk), .write_enable(1'b0), .address(LUT_address_42), .output_data(LUT_output_data_42)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_44.data") LUT_43( .clk(clk), .write_enable(1'b0), .address(LUT_address_43), .output_data(LUT_output_data_43)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_45.data") LUT_44( .clk(clk), .write_enable(1'b0), .address(LUT_address_44), .output_data(LUT_output_data_44)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_46.data") LUT_45( .clk(clk), .write_enable(1'b0), .address(LUT_address_45), .output_data(LUT_output_data_45)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_47.data") LUT_46( .clk(clk), .write_enable(1'b0), .address(LUT_address_46), .output_data(LUT_output_data_46)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_48.data") LUT_47( .clk(clk), .write_enable(1'b0), .address(LUT_address_47), .output_data(LUT_output_data_47)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_49.data") LUT_48( .clk(clk), .write_enable(1'b0), .address(LUT_address_48), .output_data(LUT_output_data_48)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_50.data") LUT_49( .clk(clk), .write_enable(1'b0), .address(LUT_address_49), .output_data(LUT_output_data_49)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_51.data") LUT_50( .clk(clk), .write_enable(1'b0), .address(LUT_address_50), .output_data(LUT_output_data_50)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_52.data") LUT_51( .clk(clk), .write_enable(1'b0), .address(LUT_address_51), .output_data(LUT_output_data_51)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_53.data") LUT_52( .clk(clk), .write_enable(1'b0), .address(LUT_address_52), .output_data(LUT_output_data_52)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_54.data") LUT_53( .clk(clk), .write_enable(1'b0), .address(LUT_address_53), .output_data(LUT_output_data_53)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_55.data") LUT_54( .clk(clk), .write_enable(1'b0), .address(LUT_address_54), .output_data(LUT_output_data_54)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_56.data") LUT_55( .clk(clk), .write_enable(1'b0), .address(LUT_address_55), .output_data(LUT_output_data_55)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_57.data") LUT_56( .clk(clk), .write_enable(1'b0), .address(LUT_address_56), .output_data(LUT_output_data_56)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_58.data") LUT_57( .clk(clk), .write_enable(1'b0), .address(LUT_address_57), .output_data(LUT_output_data_57)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_59.data") LUT_58( .clk(clk), .write_enable(1'b0), .address(LUT_address_58), .output_data(LUT_output_data_58)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_60.data") LUT_59( .clk(clk), .write_enable(1'b0), .address(LUT_address_59), .output_data(LUT_output_data_59)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_61.data") LUT_60( .clk(clk), .write_enable(1'b0), .address(LUT_address_60), .output_data(LUT_output_data_60)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_62.data") LUT_61( .clk(clk), .write_enable(1'b0), .address(LUT_address_61), .output_data(LUT_output_data_61)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_63.data") LUT_62( .clk(clk), .write_enable(1'b0), .address(LUT_address_62), .output_data(LUT_output_data_62)); 
LUT #("../../YATISH/fpgaInterfaces/ml605/preprocessed_files/1024_folding_factor_4/data/preprocessed_64.data") LUT_63( .clk(clk), .write_enable(1'b0), .address(LUT_address_63), .output_data(LUT_output_data_63)); 


endmodule

